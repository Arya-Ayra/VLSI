magic
tech scmos
timestamp 1669613447
<< nwell >>
rect -488 -508 -465 -458
rect -412 -508 -389 -458
rect -337 -508 -314 -458
rect -260 -508 -237 -458
rect -183 -508 -160 -458
rect -107 -508 -84 -458
rect -16 -508 7 -458
rect 64 -507 87 -457
rect 143 -506 166 -456
rect 219 -505 242 -455
rect 533 -504 556 -454
rect 615 -504 638 -454
rect 695 -504 718 -454
rect 824 -505 847 -455
rect 921 -505 944 -455
rect 1005 -507 1028 -457
rect -488 -564 -465 -514
rect -412 -564 -389 -514
rect -337 -564 -314 -514
rect -260 -564 -237 -514
rect -183 -564 -160 -514
rect -107 -564 -84 -514
rect -16 -564 7 -514
rect 64 -563 87 -513
rect 143 -562 166 -512
rect 219 -561 242 -511
rect 533 -560 556 -510
rect 615 -560 638 -510
rect 695 -560 718 -510
rect 824 -561 847 -511
rect 921 -561 944 -511
rect 1005 -563 1028 -513
rect 857 -639 907 -616
rect 52 -685 102 -662
rect 454 -665 504 -642
rect -467 -782 -444 -732
rect -378 -754 -355 -704
rect -139 -739 -89 -716
rect -82 -739 -32 -716
rect -3 -737 47 -714
rect 126 -715 176 -692
rect 263 -719 313 -696
rect 320 -719 370 -696
rect 399 -717 449 -694
rect 528 -695 578 -672
rect 666 -693 716 -670
rect 723 -693 773 -670
rect 802 -691 852 -668
rect 931 -669 981 -646
rect 865 -714 915 -691
rect -467 -839 -444 -789
rect -401 -817 -378 -767
rect -326 -809 -303 -759
rect 60 -760 110 -737
rect 462 -740 512 -717
rect -356 -883 -333 -833
rect -528 -965 -505 -915
rect -462 -965 -439 -915
rect -373 -966 -350 -916
rect -541 -1046 -518 -996
rect -462 -1022 -439 -972
rect -396 -1029 -373 -979
rect -321 -1021 -298 -971
rect -159 -993 -136 -943
rect -70 -965 -47 -915
rect -449 -1090 -426 -1040
rect -351 -1095 -328 -1045
rect -159 -1050 -136 -1000
rect -93 -1028 -70 -978
rect -18 -1020 5 -970
rect 174 -1012 197 -962
rect 263 -984 286 -934
rect -48 -1094 -25 -1044
rect 174 -1069 197 -1019
rect 240 -1047 263 -997
rect 315 -1039 338 -989
rect 717 -1051 740 -1001
rect 806 -1023 829 -973
rect 285 -1113 308 -1063
rect 717 -1108 740 -1058
rect 783 -1086 806 -1036
rect 858 -1078 881 -1028
rect -220 -1176 -197 -1126
rect -154 -1176 -131 -1126
rect -65 -1177 -42 -1127
rect -233 -1257 -210 -1207
rect -154 -1233 -131 -1183
rect -88 -1240 -65 -1190
rect -13 -1232 10 -1182
rect 113 -1195 136 -1145
rect 179 -1195 202 -1145
rect 268 -1196 291 -1146
rect 828 -1152 851 -1102
rect -141 -1301 -118 -1251
rect -43 -1306 -20 -1256
rect 100 -1276 123 -1226
rect 179 -1252 202 -1202
rect 245 -1259 268 -1209
rect 320 -1251 343 -1201
rect 656 -1234 679 -1184
rect 722 -1234 745 -1184
rect 811 -1235 834 -1185
rect 192 -1320 215 -1270
rect 290 -1325 313 -1275
rect 643 -1315 666 -1265
rect 722 -1291 745 -1241
rect 788 -1298 811 -1248
rect 863 -1290 886 -1240
rect 735 -1359 758 -1309
rect 833 -1364 856 -1314
rect -528 -1678 -505 -1628
rect -439 -1650 -416 -1600
rect -223 -1622 -200 -1572
rect -134 -1594 -111 -1544
rect -528 -1735 -505 -1685
rect -462 -1713 -439 -1663
rect -387 -1705 -364 -1655
rect -223 -1679 -200 -1629
rect -157 -1657 -134 -1607
rect -82 -1649 -59 -1599
rect 117 -1632 140 -1582
rect 206 -1604 229 -1554
rect 420 -1574 443 -1524
rect 509 -1546 532 -1496
rect -112 -1723 -89 -1673
rect 117 -1689 140 -1639
rect 183 -1667 206 -1617
rect 258 -1659 281 -1609
rect 420 -1631 443 -1581
rect 486 -1609 509 -1559
rect 561 -1601 584 -1551
rect 531 -1675 554 -1625
rect -417 -1779 -394 -1729
rect 228 -1733 251 -1683
rect -284 -1805 -261 -1755
rect -218 -1805 -195 -1755
rect -129 -1806 -106 -1756
rect 359 -1757 382 -1707
rect 425 -1757 448 -1707
rect 514 -1758 537 -1708
rect -589 -1861 -566 -1811
rect -523 -1861 -500 -1811
rect -434 -1862 -411 -1812
rect -602 -1942 -579 -1892
rect -523 -1918 -500 -1868
rect -457 -1925 -434 -1875
rect -382 -1917 -359 -1867
rect -297 -1886 -274 -1836
rect -218 -1862 -195 -1812
rect -152 -1869 -129 -1819
rect -77 -1861 -54 -1811
rect 56 -1815 79 -1765
rect 122 -1815 145 -1765
rect 211 -1816 234 -1766
rect -205 -1930 -182 -1880
rect -107 -1935 -84 -1885
rect 43 -1896 66 -1846
rect 122 -1872 145 -1822
rect 188 -1879 211 -1829
rect 263 -1871 286 -1821
rect 346 -1838 369 -1788
rect 425 -1814 448 -1764
rect 491 -1821 514 -1771
rect 566 -1813 589 -1763
rect 438 -1882 461 -1832
rect 536 -1887 559 -1837
rect -510 -1986 -487 -1936
rect 135 -1940 158 -1890
rect -412 -1991 -389 -1941
rect 233 -1945 256 -1895
rect 438 -2054 488 -2031
rect 247 -2108 297 -2085
rect 304 -2108 354 -2085
rect 383 -2106 433 -2083
rect 512 -2084 562 -2061
rect 446 -2129 496 -2106
<< ntransistor >>
rect -513 -473 -507 -471
rect -437 -473 -431 -471
rect -362 -473 -356 -471
rect -285 -473 -279 -471
rect -208 -473 -202 -471
rect -132 -473 -126 -471
rect -41 -473 -35 -471
rect 39 -472 45 -470
rect 118 -471 124 -469
rect 194 -470 200 -468
rect 508 -469 514 -467
rect 590 -469 596 -467
rect 670 -469 676 -467
rect 799 -470 805 -468
rect 896 -470 902 -468
rect 980 -472 986 -470
rect -513 -496 -507 -494
rect -437 -496 -431 -494
rect -362 -496 -356 -494
rect -285 -496 -279 -494
rect -208 -496 -202 -494
rect -132 -496 -126 -494
rect -41 -496 -35 -494
rect 39 -495 45 -493
rect 118 -494 124 -492
rect 194 -493 200 -491
rect 508 -492 514 -490
rect 590 -492 596 -490
rect 670 -492 676 -490
rect 799 -493 805 -491
rect 896 -493 902 -491
rect 980 -495 986 -493
rect -513 -529 -507 -527
rect -437 -529 -431 -527
rect -362 -529 -356 -527
rect -285 -529 -279 -527
rect -208 -529 -202 -527
rect -132 -529 -126 -527
rect -41 -529 -35 -527
rect 39 -528 45 -526
rect 118 -527 124 -525
rect 194 -526 200 -524
rect 508 -525 514 -523
rect 590 -525 596 -523
rect 670 -525 676 -523
rect 799 -526 805 -524
rect 896 -526 902 -524
rect 980 -528 986 -526
rect -513 -552 -507 -550
rect -437 -552 -431 -550
rect -362 -552 -356 -550
rect -285 -552 -279 -550
rect -208 -552 -202 -550
rect -132 -552 -126 -550
rect -41 -552 -35 -550
rect 39 -551 45 -549
rect 118 -550 124 -548
rect 194 -549 200 -547
rect 508 -548 514 -546
rect 590 -548 596 -546
rect 670 -548 676 -546
rect 799 -549 805 -547
rect 896 -549 902 -547
rect 980 -551 986 -549
rect 870 -664 872 -658
rect 893 -664 895 -658
rect 467 -690 469 -684
rect 490 -690 492 -684
rect 65 -710 67 -704
rect 88 -710 90 -704
rect -403 -719 -397 -717
rect -403 -742 -397 -740
rect -492 -747 -486 -745
rect 139 -740 141 -734
rect 162 -740 164 -734
rect 944 -694 946 -688
rect 967 -694 969 -688
rect 541 -720 543 -714
rect 564 -720 566 -714
rect 678 -718 680 -712
rect 701 -718 703 -712
rect 735 -718 737 -712
rect 758 -718 760 -712
rect 815 -716 817 -710
rect 838 -716 840 -710
rect 275 -744 277 -738
rect 298 -744 300 -738
rect 332 -744 334 -738
rect 355 -744 357 -738
rect 412 -742 414 -736
rect 435 -742 437 -736
rect -127 -764 -125 -758
rect -104 -764 -102 -758
rect -70 -764 -68 -758
rect -47 -764 -45 -758
rect 10 -762 12 -756
rect 33 -762 35 -756
rect -492 -770 -486 -768
rect -351 -774 -345 -772
rect 878 -739 880 -733
rect 901 -739 903 -733
rect 475 -765 477 -759
rect 498 -765 500 -759
rect -426 -782 -420 -780
rect 73 -785 75 -779
rect 96 -785 98 -779
rect -351 -797 -345 -795
rect -492 -804 -486 -802
rect -426 -805 -420 -803
rect -492 -827 -486 -825
rect -381 -848 -375 -846
rect -381 -871 -375 -869
rect -553 -930 -547 -928
rect -487 -930 -481 -928
rect -398 -931 -392 -929
rect -95 -930 -89 -928
rect -553 -953 -547 -951
rect -487 -953 -481 -951
rect 238 -949 244 -947
rect -398 -954 -392 -952
rect -95 -953 -89 -951
rect -184 -958 -178 -956
rect 238 -972 244 -970
rect 149 -977 155 -975
rect -184 -981 -178 -979
rect -487 -987 -481 -985
rect -346 -986 -340 -984
rect -43 -985 -37 -983
rect 781 -988 787 -986
rect -421 -994 -415 -992
rect -118 -993 -112 -991
rect 149 -1000 155 -998
rect 290 -1004 296 -1002
rect -566 -1011 -560 -1009
rect -487 -1010 -481 -1008
rect -346 -1009 -340 -1007
rect -43 -1008 -37 -1006
rect -184 -1015 -178 -1013
rect 215 -1012 221 -1010
rect -421 -1017 -415 -1015
rect -118 -1016 -112 -1014
rect 781 -1011 787 -1009
rect 692 -1016 698 -1014
rect 290 -1027 296 -1025
rect -566 -1034 -560 -1032
rect 149 -1034 155 -1032
rect -184 -1038 -178 -1036
rect 215 -1035 221 -1033
rect 692 -1039 698 -1037
rect 833 -1043 839 -1041
rect -474 -1055 -468 -1053
rect 758 -1051 764 -1049
rect 149 -1057 155 -1055
rect -376 -1060 -370 -1058
rect -73 -1059 -67 -1057
rect 833 -1066 839 -1064
rect -474 -1078 -468 -1076
rect 692 -1073 698 -1071
rect 260 -1078 266 -1076
rect 758 -1074 764 -1072
rect -376 -1083 -370 -1081
rect -73 -1082 -67 -1080
rect 692 -1096 698 -1094
rect 260 -1101 266 -1099
rect 803 -1117 809 -1115
rect -245 -1141 -239 -1139
rect -179 -1141 -173 -1139
rect 803 -1140 809 -1138
rect -90 -1142 -84 -1140
rect -245 -1164 -239 -1162
rect -179 -1164 -173 -1162
rect 88 -1160 94 -1158
rect 154 -1160 160 -1158
rect -90 -1165 -84 -1163
rect 243 -1161 249 -1159
rect 88 -1183 94 -1181
rect 154 -1183 160 -1181
rect 243 -1184 249 -1182
rect -179 -1198 -173 -1196
rect -38 -1197 -32 -1195
rect 631 -1199 637 -1197
rect 697 -1199 703 -1197
rect -113 -1205 -107 -1203
rect 786 -1200 792 -1198
rect 154 -1217 160 -1215
rect 295 -1216 301 -1214
rect -258 -1222 -252 -1220
rect -179 -1221 -173 -1219
rect -38 -1220 -32 -1218
rect 631 -1222 637 -1220
rect 697 -1222 703 -1220
rect 220 -1224 226 -1222
rect -113 -1228 -107 -1226
rect 786 -1223 792 -1221
rect 75 -1241 81 -1239
rect 154 -1240 160 -1238
rect 295 -1239 301 -1237
rect -258 -1245 -252 -1243
rect 220 -1247 226 -1245
rect 697 -1256 703 -1254
rect 838 -1255 844 -1253
rect 75 -1264 81 -1262
rect 763 -1263 769 -1261
rect -166 -1266 -160 -1264
rect -68 -1271 -62 -1269
rect 618 -1280 624 -1278
rect 697 -1279 703 -1277
rect 838 -1278 844 -1276
rect 167 -1285 173 -1283
rect -166 -1289 -160 -1287
rect 763 -1286 769 -1284
rect 265 -1290 271 -1288
rect -68 -1294 -62 -1292
rect 618 -1303 624 -1301
rect 167 -1308 173 -1306
rect 265 -1313 271 -1311
rect 710 -1324 716 -1322
rect 808 -1329 814 -1327
rect 710 -1347 716 -1345
rect 808 -1352 814 -1350
rect 484 -1511 490 -1509
rect 484 -1534 490 -1532
rect 395 -1539 401 -1537
rect -159 -1559 -153 -1557
rect 395 -1562 401 -1560
rect 536 -1566 542 -1564
rect 181 -1569 187 -1567
rect 461 -1574 467 -1572
rect -159 -1582 -153 -1580
rect -248 -1587 -242 -1585
rect 536 -1589 542 -1587
rect 181 -1592 187 -1590
rect 92 -1597 98 -1595
rect 395 -1596 401 -1594
rect 461 -1597 467 -1595
rect -248 -1610 -242 -1608
rect -464 -1615 -458 -1613
rect -107 -1614 -101 -1612
rect 92 -1620 98 -1618
rect -182 -1622 -176 -1620
rect 395 -1619 401 -1617
rect 233 -1624 239 -1622
rect 158 -1632 164 -1630
rect -464 -1638 -458 -1636
rect -107 -1637 -101 -1635
rect -553 -1643 -547 -1641
rect -248 -1644 -242 -1642
rect 506 -1640 512 -1638
rect -182 -1645 -176 -1643
rect 233 -1647 239 -1645
rect 92 -1654 98 -1652
rect 158 -1655 164 -1653
rect -553 -1666 -547 -1664
rect 506 -1663 512 -1661
rect -248 -1667 -242 -1665
rect -412 -1670 -406 -1668
rect -487 -1678 -481 -1676
rect 92 -1677 98 -1675
rect -137 -1688 -131 -1686
rect -412 -1693 -406 -1691
rect -553 -1700 -547 -1698
rect 203 -1698 209 -1696
rect -487 -1701 -481 -1699
rect -137 -1711 -131 -1709
rect 203 -1721 209 -1719
rect -553 -1723 -547 -1721
rect 334 -1722 340 -1720
rect 400 -1722 406 -1720
rect 489 -1723 495 -1721
rect -442 -1744 -436 -1742
rect 334 -1745 340 -1743
rect 400 -1745 406 -1743
rect 489 -1746 495 -1744
rect -442 -1767 -436 -1765
rect -309 -1770 -303 -1768
rect -243 -1770 -237 -1768
rect -154 -1771 -148 -1769
rect 31 -1780 37 -1778
rect 97 -1780 103 -1778
rect 400 -1779 406 -1777
rect 541 -1778 547 -1776
rect 186 -1781 192 -1779
rect 466 -1786 472 -1784
rect -309 -1793 -303 -1791
rect -243 -1793 -237 -1791
rect -154 -1794 -148 -1792
rect 31 -1803 37 -1801
rect 97 -1803 103 -1801
rect 186 -1804 192 -1802
rect 321 -1803 327 -1801
rect 400 -1802 406 -1800
rect 541 -1801 547 -1799
rect 466 -1809 472 -1807
rect -614 -1826 -608 -1824
rect -548 -1826 -542 -1824
rect -459 -1827 -453 -1825
rect -243 -1827 -237 -1825
rect -102 -1826 -96 -1824
rect 321 -1826 327 -1824
rect -177 -1834 -171 -1832
rect 97 -1837 103 -1835
rect 238 -1836 244 -1834
rect -614 -1849 -608 -1847
rect -548 -1849 -542 -1847
rect -459 -1850 -453 -1848
rect 163 -1844 169 -1842
rect -322 -1851 -316 -1849
rect -243 -1850 -237 -1848
rect -102 -1849 -96 -1847
rect 413 -1847 419 -1845
rect 511 -1852 517 -1850
rect -177 -1857 -171 -1855
rect 18 -1861 24 -1859
rect 97 -1860 103 -1858
rect 238 -1859 244 -1857
rect 163 -1867 169 -1865
rect 413 -1870 419 -1868
rect -322 -1874 -316 -1872
rect 511 -1875 517 -1873
rect -548 -1883 -542 -1881
rect -407 -1882 -401 -1880
rect 18 -1884 24 -1882
rect -482 -1890 -476 -1888
rect -230 -1895 -224 -1893
rect -132 -1900 -126 -1898
rect -627 -1907 -621 -1905
rect -548 -1906 -542 -1904
rect -407 -1905 -401 -1903
rect 110 -1905 116 -1903
rect 208 -1910 214 -1908
rect -482 -1913 -476 -1911
rect -230 -1918 -224 -1916
rect -132 -1923 -126 -1921
rect 110 -1928 116 -1926
rect -627 -1930 -621 -1928
rect 208 -1933 214 -1931
rect -535 -1951 -529 -1949
rect -437 -1956 -431 -1954
rect -535 -1974 -529 -1972
rect -437 -1979 -431 -1977
rect 451 -2079 453 -2073
rect 474 -2079 476 -2073
rect 525 -2109 527 -2103
rect 548 -2109 550 -2103
rect 259 -2133 261 -2127
rect 282 -2133 284 -2127
rect 316 -2133 318 -2127
rect 339 -2133 341 -2127
rect 396 -2131 398 -2125
rect 419 -2131 421 -2125
rect 459 -2154 461 -2148
rect 482 -2154 484 -2148
<< ptransistor >>
rect -481 -473 -473 -471
rect -405 -473 -397 -471
rect -330 -473 -322 -471
rect -253 -473 -245 -471
rect -176 -473 -168 -471
rect -100 -473 -92 -471
rect -9 -473 -1 -471
rect 71 -472 79 -470
rect 150 -471 158 -469
rect 226 -470 234 -468
rect 540 -469 548 -467
rect 622 -469 630 -467
rect 702 -469 710 -467
rect 831 -470 839 -468
rect 928 -470 936 -468
rect 1012 -472 1020 -470
rect -481 -496 -473 -494
rect -405 -496 -397 -494
rect -330 -496 -322 -494
rect -253 -496 -245 -494
rect -176 -496 -168 -494
rect -100 -496 -92 -494
rect -9 -496 -1 -494
rect 71 -495 79 -493
rect 150 -494 158 -492
rect 226 -493 234 -491
rect 540 -492 548 -490
rect 622 -492 630 -490
rect 702 -492 710 -490
rect 831 -493 839 -491
rect 928 -493 936 -491
rect 1012 -495 1020 -493
rect -481 -529 -473 -527
rect -405 -529 -397 -527
rect -330 -529 -322 -527
rect -253 -529 -245 -527
rect -176 -529 -168 -527
rect -100 -529 -92 -527
rect -9 -529 -1 -527
rect 71 -528 79 -526
rect 150 -527 158 -525
rect 226 -526 234 -524
rect 540 -525 548 -523
rect 622 -525 630 -523
rect 702 -525 710 -523
rect 831 -526 839 -524
rect 928 -526 936 -524
rect 1012 -528 1020 -526
rect -481 -552 -473 -550
rect -405 -552 -397 -550
rect -330 -552 -322 -550
rect -253 -552 -245 -550
rect -176 -552 -168 -550
rect -100 -552 -92 -550
rect -9 -552 -1 -550
rect 71 -551 79 -549
rect 150 -550 158 -548
rect 226 -549 234 -547
rect 540 -548 548 -546
rect 622 -548 630 -546
rect 702 -548 710 -546
rect 831 -549 839 -547
rect 928 -549 936 -547
rect 1012 -551 1020 -549
rect 870 -632 872 -624
rect 893 -632 895 -624
rect 467 -658 469 -650
rect 490 -658 492 -650
rect 65 -678 67 -670
rect 88 -678 90 -670
rect 944 -662 946 -654
rect 967 -662 969 -654
rect 541 -688 543 -680
rect 564 -688 566 -680
rect 678 -686 680 -678
rect 701 -686 703 -678
rect 735 -686 737 -678
rect 758 -686 760 -678
rect 815 -684 817 -676
rect 838 -684 840 -676
rect 139 -708 141 -700
rect 162 -708 164 -700
rect -371 -719 -363 -717
rect -127 -732 -125 -724
rect -104 -732 -102 -724
rect -70 -732 -68 -724
rect -47 -732 -45 -724
rect 10 -730 12 -722
rect 33 -730 35 -722
rect -371 -742 -363 -740
rect -460 -747 -452 -745
rect 275 -712 277 -704
rect 298 -712 300 -704
rect 332 -712 334 -704
rect 355 -712 357 -704
rect 412 -710 414 -702
rect 435 -710 437 -702
rect 878 -707 880 -699
rect 901 -707 903 -699
rect 475 -733 477 -725
rect 498 -733 500 -725
rect 73 -753 75 -745
rect 96 -753 98 -745
rect -460 -770 -452 -768
rect -319 -774 -311 -772
rect -394 -782 -386 -780
rect -319 -797 -311 -795
rect -460 -804 -452 -802
rect -394 -805 -386 -803
rect -460 -827 -452 -825
rect -349 -848 -341 -846
rect -349 -871 -341 -869
rect -521 -930 -513 -928
rect -455 -930 -447 -928
rect -366 -931 -358 -929
rect -63 -930 -55 -928
rect -521 -953 -513 -951
rect -455 -953 -447 -951
rect 270 -949 278 -947
rect -366 -954 -358 -952
rect -63 -953 -55 -951
rect -152 -958 -144 -956
rect 270 -972 278 -970
rect 181 -977 189 -975
rect -152 -981 -144 -979
rect -455 -987 -447 -985
rect -314 -986 -306 -984
rect -11 -985 -3 -983
rect 813 -988 821 -986
rect -389 -994 -381 -992
rect -86 -993 -78 -991
rect 181 -1000 189 -998
rect 322 -1004 330 -1002
rect -534 -1011 -526 -1009
rect -455 -1010 -447 -1008
rect -314 -1009 -306 -1007
rect -11 -1008 -3 -1006
rect -152 -1015 -144 -1013
rect 247 -1012 255 -1010
rect -389 -1017 -381 -1015
rect -86 -1016 -78 -1014
rect 813 -1011 821 -1009
rect 724 -1016 732 -1014
rect 322 -1027 330 -1025
rect -534 -1034 -526 -1032
rect 181 -1034 189 -1032
rect -152 -1038 -144 -1036
rect 247 -1035 255 -1033
rect 724 -1039 732 -1037
rect 865 -1043 873 -1041
rect -442 -1055 -434 -1053
rect 790 -1051 798 -1049
rect 181 -1057 189 -1055
rect -344 -1060 -336 -1058
rect -41 -1059 -33 -1057
rect 865 -1066 873 -1064
rect -442 -1078 -434 -1076
rect 724 -1073 732 -1071
rect 292 -1078 300 -1076
rect 790 -1074 798 -1072
rect -344 -1083 -336 -1081
rect -41 -1082 -33 -1080
rect 724 -1096 732 -1094
rect 292 -1101 300 -1099
rect 835 -1117 843 -1115
rect -213 -1141 -205 -1139
rect -147 -1141 -139 -1139
rect 835 -1140 843 -1138
rect -58 -1142 -50 -1140
rect -213 -1164 -205 -1162
rect -147 -1164 -139 -1162
rect 120 -1160 128 -1158
rect 186 -1160 194 -1158
rect -58 -1165 -50 -1163
rect 275 -1161 283 -1159
rect 120 -1183 128 -1181
rect 186 -1183 194 -1181
rect 275 -1184 283 -1182
rect -147 -1198 -139 -1196
rect -6 -1197 2 -1195
rect 663 -1199 671 -1197
rect 729 -1199 737 -1197
rect -81 -1205 -73 -1203
rect 818 -1200 826 -1198
rect 186 -1217 194 -1215
rect 327 -1216 335 -1214
rect -226 -1222 -218 -1220
rect -147 -1221 -139 -1219
rect -6 -1220 2 -1218
rect 663 -1222 671 -1220
rect 729 -1222 737 -1220
rect 252 -1224 260 -1222
rect -81 -1228 -73 -1226
rect 818 -1223 826 -1221
rect 107 -1241 115 -1239
rect 186 -1240 194 -1238
rect 327 -1239 335 -1237
rect -226 -1245 -218 -1243
rect 252 -1247 260 -1245
rect 729 -1256 737 -1254
rect 870 -1255 878 -1253
rect 107 -1264 115 -1262
rect 795 -1263 803 -1261
rect -134 -1266 -126 -1264
rect -36 -1271 -28 -1269
rect 650 -1280 658 -1278
rect 729 -1279 737 -1277
rect 870 -1278 878 -1276
rect 199 -1285 207 -1283
rect -134 -1289 -126 -1287
rect 795 -1286 803 -1284
rect 297 -1290 305 -1288
rect -36 -1294 -28 -1292
rect 650 -1303 658 -1301
rect 199 -1308 207 -1306
rect 297 -1313 305 -1311
rect 742 -1324 750 -1322
rect 840 -1329 848 -1327
rect 742 -1347 750 -1345
rect 840 -1352 848 -1350
rect 516 -1511 524 -1509
rect 516 -1534 524 -1532
rect 427 -1539 435 -1537
rect -127 -1559 -119 -1557
rect 427 -1562 435 -1560
rect 568 -1566 576 -1564
rect 213 -1569 221 -1567
rect 493 -1574 501 -1572
rect -127 -1582 -119 -1580
rect -216 -1587 -208 -1585
rect 568 -1589 576 -1587
rect 213 -1592 221 -1590
rect 124 -1597 132 -1595
rect 427 -1596 435 -1594
rect 493 -1597 501 -1595
rect -216 -1610 -208 -1608
rect -432 -1615 -424 -1613
rect -75 -1614 -67 -1612
rect 124 -1620 132 -1618
rect -150 -1622 -142 -1620
rect 427 -1619 435 -1617
rect 265 -1624 273 -1622
rect 190 -1632 198 -1630
rect -432 -1638 -424 -1636
rect -75 -1637 -67 -1635
rect -521 -1643 -513 -1641
rect -216 -1644 -208 -1642
rect 538 -1640 546 -1638
rect -150 -1645 -142 -1643
rect 265 -1647 273 -1645
rect 124 -1654 132 -1652
rect 190 -1655 198 -1653
rect -521 -1666 -513 -1664
rect 538 -1663 546 -1661
rect -216 -1667 -208 -1665
rect -380 -1670 -372 -1668
rect -455 -1678 -447 -1676
rect 124 -1677 132 -1675
rect -105 -1688 -97 -1686
rect -380 -1693 -372 -1691
rect -521 -1700 -513 -1698
rect 235 -1698 243 -1696
rect -455 -1701 -447 -1699
rect -105 -1711 -97 -1709
rect 235 -1721 243 -1719
rect -521 -1723 -513 -1721
rect 366 -1722 374 -1720
rect 432 -1722 440 -1720
rect 521 -1723 529 -1721
rect -410 -1744 -402 -1742
rect 366 -1745 374 -1743
rect 432 -1745 440 -1743
rect 521 -1746 529 -1744
rect -410 -1767 -402 -1765
rect -277 -1770 -269 -1768
rect -211 -1770 -203 -1768
rect -122 -1771 -114 -1769
rect 63 -1780 71 -1778
rect 129 -1780 137 -1778
rect 432 -1779 440 -1777
rect 573 -1778 581 -1776
rect 218 -1781 226 -1779
rect 498 -1786 506 -1784
rect -277 -1793 -269 -1791
rect -211 -1793 -203 -1791
rect -122 -1794 -114 -1792
rect 63 -1803 71 -1801
rect 129 -1803 137 -1801
rect 218 -1804 226 -1802
rect 353 -1803 361 -1801
rect 432 -1802 440 -1800
rect 573 -1801 581 -1799
rect 498 -1809 506 -1807
rect -582 -1826 -574 -1824
rect -516 -1826 -508 -1824
rect -427 -1827 -419 -1825
rect -211 -1827 -203 -1825
rect -70 -1826 -62 -1824
rect 353 -1826 361 -1824
rect -145 -1834 -137 -1832
rect 129 -1837 137 -1835
rect 270 -1836 278 -1834
rect -582 -1849 -574 -1847
rect -516 -1849 -508 -1847
rect -427 -1850 -419 -1848
rect 195 -1844 203 -1842
rect -290 -1851 -282 -1849
rect -211 -1850 -203 -1848
rect -70 -1849 -62 -1847
rect 445 -1847 453 -1845
rect 543 -1852 551 -1850
rect -145 -1857 -137 -1855
rect 50 -1861 58 -1859
rect 129 -1860 137 -1858
rect 270 -1859 278 -1857
rect 195 -1867 203 -1865
rect 445 -1870 453 -1868
rect -290 -1874 -282 -1872
rect 543 -1875 551 -1873
rect -516 -1883 -508 -1881
rect -375 -1882 -367 -1880
rect 50 -1884 58 -1882
rect -450 -1890 -442 -1888
rect -198 -1895 -190 -1893
rect -100 -1900 -92 -1898
rect -595 -1907 -587 -1905
rect -516 -1906 -508 -1904
rect -375 -1905 -367 -1903
rect 142 -1905 150 -1903
rect 240 -1910 248 -1908
rect -450 -1913 -442 -1911
rect -198 -1918 -190 -1916
rect -100 -1923 -92 -1921
rect 142 -1928 150 -1926
rect -595 -1930 -587 -1928
rect 240 -1933 248 -1931
rect -503 -1951 -495 -1949
rect -405 -1956 -397 -1954
rect -503 -1974 -495 -1972
rect -405 -1979 -397 -1977
rect 451 -2047 453 -2039
rect 474 -2047 476 -2039
rect 525 -2077 527 -2069
rect 548 -2077 550 -2069
rect 259 -2101 261 -2093
rect 282 -2101 284 -2093
rect 316 -2101 318 -2093
rect 339 -2101 341 -2093
rect 396 -2099 398 -2091
rect 419 -2099 421 -2091
rect 459 -2122 461 -2114
rect 482 -2122 484 -2114
<< ndiffusion >>
rect -513 -471 -507 -470
rect -437 -471 -431 -470
rect -362 -471 -356 -470
rect -285 -471 -279 -470
rect -208 -471 -202 -470
rect -132 -471 -126 -470
rect -41 -471 -35 -470
rect 39 -470 45 -469
rect 118 -469 124 -468
rect 194 -468 200 -467
rect 508 -467 514 -466
rect 590 -467 596 -466
rect 670 -467 676 -466
rect 799 -468 805 -467
rect 896 -468 902 -467
rect 508 -470 514 -469
rect 194 -471 200 -470
rect 118 -472 124 -471
rect 39 -473 45 -472
rect -513 -474 -507 -473
rect -437 -474 -431 -473
rect -362 -474 -356 -473
rect -285 -474 -279 -473
rect -208 -474 -202 -473
rect -132 -474 -126 -473
rect -41 -474 -35 -473
rect 590 -470 596 -469
rect 670 -470 676 -469
rect 980 -470 986 -469
rect 799 -471 805 -470
rect 896 -471 902 -470
rect 980 -473 986 -472
rect -513 -494 -507 -493
rect -437 -494 -431 -493
rect -362 -494 -356 -493
rect -285 -494 -279 -493
rect -208 -494 -202 -493
rect -132 -494 -126 -493
rect -41 -494 -35 -493
rect 39 -493 45 -492
rect 118 -492 124 -491
rect 194 -491 200 -490
rect 508 -490 514 -489
rect 590 -490 596 -489
rect 670 -490 676 -489
rect 799 -491 805 -490
rect 896 -491 902 -490
rect 508 -493 514 -492
rect 194 -494 200 -493
rect 118 -495 124 -494
rect 39 -496 45 -495
rect -513 -497 -507 -496
rect -437 -497 -431 -496
rect -362 -497 -356 -496
rect -285 -497 -279 -496
rect -208 -497 -202 -496
rect -132 -497 -126 -496
rect -41 -497 -35 -496
rect 590 -493 596 -492
rect 670 -493 676 -492
rect 980 -493 986 -492
rect 799 -494 805 -493
rect 896 -494 902 -493
rect 980 -496 986 -495
rect -513 -527 -507 -526
rect -437 -527 -431 -526
rect -362 -527 -356 -526
rect -285 -527 -279 -526
rect -208 -527 -202 -526
rect -132 -527 -126 -526
rect -41 -527 -35 -526
rect 39 -526 45 -525
rect 118 -525 124 -524
rect 194 -524 200 -523
rect 508 -523 514 -522
rect 590 -523 596 -522
rect 670 -523 676 -522
rect 799 -524 805 -523
rect 896 -524 902 -523
rect 508 -526 514 -525
rect 194 -527 200 -526
rect 118 -528 124 -527
rect 39 -529 45 -528
rect -513 -530 -507 -529
rect -437 -530 -431 -529
rect -362 -530 -356 -529
rect -285 -530 -279 -529
rect -208 -530 -202 -529
rect -132 -530 -126 -529
rect -41 -530 -35 -529
rect 590 -526 596 -525
rect 670 -526 676 -525
rect 980 -526 986 -525
rect 799 -527 805 -526
rect 896 -527 902 -526
rect 980 -529 986 -528
rect -513 -550 -507 -549
rect -437 -550 -431 -549
rect -362 -550 -356 -549
rect -285 -550 -279 -549
rect -208 -550 -202 -549
rect -132 -550 -126 -549
rect -41 -550 -35 -549
rect 39 -549 45 -548
rect 118 -548 124 -547
rect 194 -547 200 -546
rect 508 -546 514 -545
rect 590 -546 596 -545
rect 670 -546 676 -545
rect 799 -547 805 -546
rect 896 -547 902 -546
rect 508 -549 514 -548
rect 194 -550 200 -549
rect 118 -551 124 -550
rect 39 -552 45 -551
rect -513 -553 -507 -552
rect -437 -553 -431 -552
rect -362 -553 -356 -552
rect -285 -553 -279 -552
rect -208 -553 -202 -552
rect -132 -553 -126 -552
rect -41 -553 -35 -552
rect 590 -549 596 -548
rect 670 -549 676 -548
rect 980 -549 986 -548
rect 799 -550 805 -549
rect 896 -550 902 -549
rect 980 -552 986 -551
rect 869 -664 870 -658
rect 872 -664 873 -658
rect 892 -664 893 -658
rect 895 -664 896 -658
rect 466 -690 467 -684
rect 469 -690 470 -684
rect 489 -690 490 -684
rect 492 -690 493 -684
rect 64 -710 65 -704
rect 67 -710 68 -704
rect 87 -710 88 -704
rect 90 -710 91 -704
rect -403 -717 -397 -716
rect -403 -720 -397 -719
rect -403 -740 -397 -739
rect -492 -745 -486 -744
rect -403 -743 -397 -742
rect -492 -748 -486 -747
rect 138 -740 139 -734
rect 141 -740 142 -734
rect 161 -740 162 -734
rect 164 -740 165 -734
rect 943 -694 944 -688
rect 946 -694 947 -688
rect 966 -694 967 -688
rect 969 -694 970 -688
rect 540 -720 541 -714
rect 543 -720 544 -714
rect 563 -720 564 -714
rect 566 -720 567 -714
rect 677 -718 678 -712
rect 680 -718 681 -712
rect 700 -718 701 -712
rect 703 -718 704 -712
rect 734 -718 735 -712
rect 737 -718 738 -712
rect 757 -718 758 -712
rect 760 -718 761 -712
rect 814 -716 815 -710
rect 817 -716 818 -710
rect 837 -716 838 -710
rect 840 -716 841 -710
rect 274 -744 275 -738
rect 277 -744 278 -738
rect 297 -744 298 -738
rect 300 -744 301 -738
rect 331 -744 332 -738
rect 334 -744 335 -738
rect 354 -744 355 -738
rect 357 -744 358 -738
rect 411 -742 412 -736
rect 414 -742 415 -736
rect 434 -742 435 -736
rect 437 -742 438 -736
rect -492 -768 -486 -767
rect -128 -764 -127 -758
rect -125 -764 -124 -758
rect -105 -764 -104 -758
rect -102 -764 -101 -758
rect -71 -764 -70 -758
rect -68 -764 -67 -758
rect -48 -764 -47 -758
rect -45 -764 -44 -758
rect 9 -762 10 -756
rect 12 -762 13 -756
rect 32 -762 33 -756
rect 35 -762 36 -756
rect -492 -771 -486 -770
rect -351 -772 -345 -771
rect -351 -775 -345 -774
rect -426 -780 -420 -779
rect 877 -739 878 -733
rect 880 -739 881 -733
rect 900 -739 901 -733
rect 903 -739 904 -733
rect 474 -765 475 -759
rect 477 -765 478 -759
rect 497 -765 498 -759
rect 500 -765 501 -759
rect -426 -783 -420 -782
rect 72 -785 73 -779
rect 75 -785 76 -779
rect 95 -785 96 -779
rect 98 -785 99 -779
rect -351 -795 -345 -794
rect -492 -802 -486 -801
rect -351 -798 -345 -797
rect -426 -803 -420 -802
rect -492 -805 -486 -804
rect -426 -806 -420 -805
rect -492 -825 -486 -824
rect -492 -828 -486 -827
rect -381 -846 -375 -845
rect -381 -849 -375 -848
rect -381 -869 -375 -868
rect -381 -872 -375 -871
rect -553 -928 -547 -927
rect -487 -928 -481 -927
rect -398 -929 -392 -928
rect -95 -928 -89 -927
rect -553 -931 -547 -930
rect -487 -931 -481 -930
rect -95 -931 -89 -930
rect -398 -932 -392 -931
rect -553 -951 -547 -950
rect -487 -951 -481 -950
rect -398 -952 -392 -951
rect -95 -951 -89 -950
rect 238 -947 244 -946
rect 238 -950 244 -949
rect -553 -954 -547 -953
rect -487 -954 -481 -953
rect -398 -955 -392 -954
rect -184 -956 -178 -955
rect -95 -954 -89 -953
rect -184 -959 -178 -958
rect 238 -970 244 -969
rect -184 -979 -178 -978
rect 149 -975 155 -974
rect 238 -973 244 -972
rect 149 -978 155 -977
rect -487 -985 -481 -984
rect -346 -984 -340 -983
rect -184 -982 -178 -981
rect -43 -983 -37 -982
rect -43 -986 -37 -985
rect -346 -987 -340 -986
rect -487 -988 -481 -987
rect -421 -992 -415 -991
rect -118 -991 -112 -990
rect 781 -986 787 -985
rect 781 -989 787 -988
rect -118 -994 -112 -993
rect -421 -995 -415 -994
rect 149 -998 155 -997
rect 149 -1001 155 -1000
rect -566 -1009 -560 -1008
rect -487 -1008 -481 -1007
rect -346 -1007 -340 -1006
rect -43 -1006 -37 -1005
rect 290 -1002 296 -1001
rect 290 -1005 296 -1004
rect -346 -1010 -340 -1009
rect -487 -1011 -481 -1010
rect -566 -1012 -560 -1011
rect -421 -1015 -415 -1014
rect -184 -1013 -178 -1012
rect -43 -1009 -37 -1008
rect -118 -1014 -112 -1013
rect 215 -1010 221 -1009
rect 781 -1009 787 -1008
rect 215 -1013 221 -1012
rect -184 -1016 -178 -1015
rect -421 -1018 -415 -1017
rect -118 -1017 -112 -1016
rect 692 -1014 698 -1013
rect 781 -1012 787 -1011
rect 692 -1017 698 -1016
rect 290 -1025 296 -1024
rect -566 -1032 -560 -1031
rect -566 -1035 -560 -1034
rect -184 -1036 -178 -1035
rect 149 -1032 155 -1031
rect 290 -1028 296 -1027
rect 215 -1033 221 -1032
rect 149 -1035 155 -1034
rect -184 -1039 -178 -1038
rect 215 -1036 221 -1035
rect 692 -1037 698 -1036
rect 692 -1040 698 -1039
rect 833 -1041 839 -1040
rect 833 -1044 839 -1043
rect -474 -1053 -468 -1052
rect 758 -1049 764 -1048
rect -474 -1056 -468 -1055
rect -376 -1058 -370 -1057
rect -73 -1057 -67 -1056
rect 149 -1055 155 -1054
rect 758 -1052 764 -1051
rect 149 -1058 155 -1057
rect -73 -1060 -67 -1059
rect -376 -1061 -370 -1060
rect 833 -1064 839 -1063
rect 692 -1071 698 -1070
rect 833 -1067 839 -1066
rect -474 -1076 -468 -1075
rect -474 -1079 -468 -1078
rect -376 -1081 -370 -1080
rect -73 -1080 -67 -1079
rect 260 -1076 266 -1075
rect 758 -1072 764 -1071
rect 692 -1074 698 -1073
rect 758 -1075 764 -1074
rect 260 -1079 266 -1078
rect -73 -1083 -67 -1082
rect -376 -1084 -370 -1083
rect 692 -1094 698 -1093
rect 260 -1099 266 -1098
rect 692 -1097 698 -1096
rect 260 -1102 266 -1101
rect 803 -1115 809 -1114
rect 803 -1118 809 -1117
rect -245 -1139 -239 -1138
rect -179 -1139 -173 -1138
rect -90 -1140 -84 -1139
rect 803 -1138 809 -1137
rect -245 -1142 -239 -1141
rect -179 -1142 -173 -1141
rect 803 -1141 809 -1140
rect -90 -1143 -84 -1142
rect -245 -1162 -239 -1161
rect -179 -1162 -173 -1161
rect 88 -1158 94 -1157
rect 154 -1158 160 -1157
rect -90 -1163 -84 -1162
rect 243 -1159 249 -1158
rect 88 -1161 94 -1160
rect -245 -1165 -239 -1164
rect -179 -1165 -173 -1164
rect 154 -1161 160 -1160
rect 243 -1162 249 -1161
rect -90 -1166 -84 -1165
rect 88 -1181 94 -1180
rect 154 -1181 160 -1180
rect 243 -1182 249 -1181
rect 88 -1184 94 -1183
rect 154 -1184 160 -1183
rect 243 -1185 249 -1184
rect -179 -1196 -173 -1195
rect -38 -1195 -32 -1194
rect 631 -1197 637 -1196
rect 697 -1197 703 -1196
rect -38 -1198 -32 -1197
rect -179 -1199 -173 -1198
rect -113 -1203 -107 -1202
rect 786 -1198 792 -1197
rect 631 -1200 637 -1199
rect 697 -1200 703 -1199
rect 786 -1201 792 -1200
rect -113 -1206 -107 -1205
rect -258 -1220 -252 -1219
rect -179 -1219 -173 -1218
rect -38 -1218 -32 -1217
rect 154 -1215 160 -1214
rect 295 -1214 301 -1213
rect 295 -1217 301 -1216
rect 154 -1218 160 -1217
rect -38 -1221 -32 -1220
rect -179 -1222 -173 -1221
rect -258 -1223 -252 -1222
rect -113 -1226 -107 -1225
rect 220 -1222 226 -1221
rect 631 -1220 637 -1219
rect 697 -1220 703 -1219
rect 786 -1221 792 -1220
rect 631 -1223 637 -1222
rect 220 -1225 226 -1224
rect -113 -1229 -107 -1228
rect 697 -1223 703 -1222
rect 786 -1224 792 -1223
rect -258 -1243 -252 -1242
rect 75 -1239 81 -1238
rect 154 -1238 160 -1237
rect 295 -1237 301 -1236
rect 295 -1240 301 -1239
rect 154 -1241 160 -1240
rect 75 -1242 81 -1241
rect -258 -1246 -252 -1245
rect 220 -1245 226 -1244
rect 220 -1248 226 -1247
rect 697 -1254 703 -1253
rect 838 -1253 844 -1252
rect 838 -1256 844 -1255
rect 697 -1257 703 -1256
rect -166 -1264 -160 -1263
rect 75 -1262 81 -1261
rect 763 -1261 769 -1260
rect 763 -1264 769 -1263
rect -166 -1267 -160 -1266
rect -68 -1269 -62 -1268
rect 75 -1265 81 -1264
rect -68 -1272 -62 -1271
rect 618 -1278 624 -1277
rect 697 -1277 703 -1276
rect 838 -1276 844 -1275
rect -166 -1287 -160 -1286
rect 167 -1283 173 -1282
rect 838 -1279 844 -1278
rect 697 -1280 703 -1279
rect 618 -1281 624 -1280
rect 167 -1286 173 -1285
rect -166 -1290 -160 -1289
rect -68 -1292 -62 -1291
rect 265 -1288 271 -1287
rect 763 -1284 769 -1283
rect 763 -1287 769 -1286
rect 265 -1291 271 -1290
rect -68 -1295 -62 -1294
rect 618 -1301 624 -1300
rect 167 -1306 173 -1305
rect 618 -1304 624 -1303
rect 167 -1309 173 -1308
rect 265 -1311 271 -1310
rect 265 -1314 271 -1313
rect 710 -1322 716 -1321
rect 710 -1325 716 -1324
rect 808 -1327 814 -1326
rect 808 -1330 814 -1329
rect 710 -1345 716 -1344
rect 710 -1348 716 -1347
rect 808 -1350 814 -1349
rect 808 -1353 814 -1352
rect 484 -1509 490 -1508
rect 484 -1512 490 -1511
rect 484 -1532 490 -1531
rect 395 -1537 401 -1536
rect 484 -1535 490 -1534
rect 395 -1540 401 -1539
rect -159 -1557 -153 -1556
rect -159 -1560 -153 -1559
rect 395 -1560 401 -1559
rect 181 -1567 187 -1566
rect 395 -1563 401 -1562
rect 536 -1564 542 -1563
rect 536 -1567 542 -1566
rect 181 -1570 187 -1569
rect 461 -1572 467 -1571
rect 461 -1575 467 -1574
rect -159 -1580 -153 -1579
rect -248 -1585 -242 -1584
rect -159 -1583 -153 -1582
rect -248 -1588 -242 -1587
rect 181 -1590 187 -1589
rect 536 -1587 542 -1586
rect 92 -1595 98 -1594
rect 181 -1593 187 -1592
rect 395 -1594 401 -1593
rect 536 -1590 542 -1589
rect 461 -1595 467 -1594
rect 395 -1597 401 -1596
rect 92 -1598 98 -1597
rect 461 -1598 467 -1597
rect -248 -1608 -242 -1607
rect -464 -1613 -458 -1612
rect -248 -1611 -242 -1610
rect -107 -1612 -101 -1611
rect -107 -1615 -101 -1614
rect -464 -1616 -458 -1615
rect -182 -1620 -176 -1619
rect 92 -1618 98 -1617
rect 395 -1617 401 -1616
rect 92 -1621 98 -1620
rect -182 -1623 -176 -1622
rect 233 -1622 239 -1621
rect 395 -1620 401 -1619
rect 233 -1625 239 -1624
rect 158 -1630 164 -1629
rect -464 -1636 -458 -1635
rect -107 -1635 -101 -1634
rect 158 -1633 164 -1632
rect -553 -1641 -547 -1640
rect -464 -1639 -458 -1638
rect -248 -1642 -242 -1641
rect -107 -1638 -101 -1637
rect -553 -1644 -547 -1643
rect -182 -1643 -176 -1642
rect 506 -1638 512 -1637
rect -248 -1645 -242 -1644
rect 233 -1645 239 -1644
rect 506 -1641 512 -1640
rect -182 -1646 -176 -1645
rect 92 -1652 98 -1651
rect 233 -1648 239 -1647
rect 158 -1653 164 -1652
rect 92 -1655 98 -1654
rect 158 -1656 164 -1655
rect -553 -1664 -547 -1663
rect -553 -1667 -547 -1666
rect -412 -1668 -406 -1667
rect -248 -1665 -242 -1664
rect 506 -1661 512 -1660
rect 506 -1664 512 -1663
rect -248 -1668 -242 -1667
rect -412 -1671 -406 -1670
rect -487 -1676 -481 -1675
rect 92 -1675 98 -1674
rect 92 -1678 98 -1677
rect -487 -1679 -481 -1678
rect -137 -1686 -131 -1685
rect -412 -1691 -406 -1690
rect -137 -1689 -131 -1688
rect -553 -1698 -547 -1697
rect -412 -1694 -406 -1693
rect -487 -1699 -481 -1698
rect 203 -1696 209 -1695
rect 203 -1699 209 -1698
rect -553 -1701 -547 -1700
rect -487 -1702 -481 -1701
rect -137 -1709 -131 -1708
rect -137 -1712 -131 -1711
rect -553 -1721 -547 -1720
rect 203 -1719 209 -1718
rect 334 -1720 340 -1719
rect 400 -1720 406 -1719
rect 203 -1722 209 -1721
rect -553 -1724 -547 -1723
rect 489 -1721 495 -1720
rect 334 -1723 340 -1722
rect 400 -1723 406 -1722
rect 489 -1724 495 -1723
rect -442 -1742 -436 -1741
rect 334 -1743 340 -1742
rect 400 -1743 406 -1742
rect -442 -1745 -436 -1744
rect 489 -1744 495 -1743
rect 334 -1746 340 -1745
rect 400 -1746 406 -1745
rect 489 -1747 495 -1746
rect -442 -1765 -436 -1764
rect -442 -1768 -436 -1767
rect -309 -1768 -303 -1767
rect -243 -1768 -237 -1767
rect -154 -1769 -148 -1768
rect -309 -1771 -303 -1770
rect -243 -1771 -237 -1770
rect -154 -1772 -148 -1771
rect 31 -1778 37 -1777
rect 97 -1778 103 -1777
rect 186 -1779 192 -1778
rect 400 -1777 406 -1776
rect 541 -1776 547 -1775
rect 541 -1779 547 -1778
rect 31 -1781 37 -1780
rect 97 -1781 103 -1780
rect 400 -1780 406 -1779
rect 186 -1782 192 -1781
rect 466 -1784 472 -1783
rect -309 -1791 -303 -1790
rect -243 -1791 -237 -1790
rect 466 -1787 472 -1786
rect -154 -1792 -148 -1791
rect -309 -1794 -303 -1793
rect -243 -1794 -237 -1793
rect -154 -1795 -148 -1794
rect 31 -1801 37 -1800
rect 97 -1801 103 -1800
rect 186 -1802 192 -1801
rect 321 -1801 327 -1800
rect 400 -1800 406 -1799
rect 541 -1799 547 -1798
rect 31 -1804 37 -1803
rect 97 -1804 103 -1803
rect 541 -1802 547 -1801
rect 400 -1803 406 -1802
rect 321 -1804 327 -1803
rect 186 -1805 192 -1804
rect 466 -1807 472 -1806
rect 466 -1810 472 -1809
rect -614 -1824 -608 -1823
rect -548 -1824 -542 -1823
rect -459 -1825 -453 -1824
rect -243 -1825 -237 -1824
rect -102 -1824 -96 -1823
rect 321 -1824 327 -1823
rect -614 -1827 -608 -1826
rect -548 -1827 -542 -1826
rect -102 -1827 -96 -1826
rect -459 -1828 -453 -1827
rect -243 -1828 -237 -1827
rect -177 -1832 -171 -1831
rect 321 -1827 327 -1826
rect -177 -1835 -171 -1834
rect 97 -1835 103 -1834
rect 238 -1834 244 -1833
rect 238 -1837 244 -1836
rect 97 -1838 103 -1837
rect 163 -1842 169 -1841
rect -614 -1847 -608 -1846
rect -548 -1847 -542 -1846
rect -459 -1848 -453 -1847
rect -614 -1850 -608 -1849
rect -548 -1850 -542 -1849
rect -322 -1849 -316 -1848
rect -243 -1848 -237 -1847
rect -102 -1847 -96 -1846
rect 163 -1845 169 -1844
rect -459 -1851 -453 -1850
rect 413 -1845 419 -1844
rect 413 -1848 419 -1847
rect -102 -1850 -96 -1849
rect -243 -1851 -237 -1850
rect -322 -1852 -316 -1851
rect -177 -1855 -171 -1854
rect 511 -1850 517 -1849
rect -177 -1858 -171 -1857
rect 18 -1859 24 -1858
rect 97 -1858 103 -1857
rect 238 -1857 244 -1856
rect 511 -1853 517 -1852
rect 238 -1860 244 -1859
rect 97 -1861 103 -1860
rect 18 -1862 24 -1861
rect 163 -1865 169 -1864
rect -322 -1872 -316 -1871
rect 163 -1868 169 -1867
rect 413 -1868 419 -1867
rect 413 -1871 419 -1870
rect -322 -1875 -316 -1874
rect -548 -1881 -542 -1880
rect -407 -1880 -401 -1879
rect 511 -1873 517 -1872
rect 511 -1876 517 -1875
rect 18 -1882 24 -1881
rect -407 -1883 -401 -1882
rect -548 -1884 -542 -1883
rect -482 -1888 -476 -1887
rect 18 -1885 24 -1884
rect -482 -1891 -476 -1890
rect -230 -1893 -224 -1892
rect -230 -1896 -224 -1895
rect -627 -1905 -621 -1904
rect -548 -1904 -542 -1903
rect -407 -1903 -401 -1902
rect -132 -1898 -126 -1897
rect -132 -1901 -126 -1900
rect 110 -1903 116 -1902
rect -407 -1906 -401 -1905
rect -548 -1907 -542 -1906
rect -627 -1908 -621 -1907
rect -482 -1911 -476 -1910
rect 110 -1906 116 -1905
rect 208 -1908 214 -1907
rect 208 -1911 214 -1910
rect -482 -1914 -476 -1913
rect -230 -1916 -224 -1915
rect -230 -1919 -224 -1918
rect -132 -1921 -126 -1920
rect -627 -1928 -621 -1927
rect -132 -1924 -126 -1923
rect 110 -1926 116 -1925
rect 110 -1929 116 -1928
rect -627 -1931 -621 -1930
rect 208 -1931 214 -1930
rect 208 -1934 214 -1933
rect -535 -1949 -529 -1948
rect -535 -1952 -529 -1951
rect -437 -1954 -431 -1953
rect -437 -1957 -431 -1956
rect -535 -1972 -529 -1971
rect -535 -1975 -529 -1974
rect -437 -1977 -431 -1976
rect -437 -1980 -431 -1979
rect 450 -2079 451 -2073
rect 453 -2079 454 -2073
rect 473 -2079 474 -2073
rect 476 -2079 477 -2073
rect 524 -2109 525 -2103
rect 527 -2109 528 -2103
rect 547 -2109 548 -2103
rect 550 -2109 551 -2103
rect 258 -2133 259 -2127
rect 261 -2133 262 -2127
rect 281 -2133 282 -2127
rect 284 -2133 285 -2127
rect 315 -2133 316 -2127
rect 318 -2133 319 -2127
rect 338 -2133 339 -2127
rect 341 -2133 342 -2127
rect 395 -2131 396 -2125
rect 398 -2131 399 -2125
rect 418 -2131 419 -2125
rect 421 -2131 422 -2125
rect 458 -2154 459 -2148
rect 461 -2154 462 -2148
rect 481 -2154 482 -2148
rect 484 -2154 485 -2148
<< pdiffusion >>
rect -481 -471 -473 -470
rect -405 -471 -397 -470
rect -330 -471 -322 -470
rect -253 -471 -245 -470
rect -176 -471 -168 -470
rect -100 -471 -92 -470
rect 540 -467 548 -466
rect 622 -467 630 -466
rect 702 -467 710 -466
rect 226 -468 234 -467
rect 150 -469 158 -468
rect 71 -470 79 -469
rect -9 -471 -1 -470
rect 831 -468 839 -467
rect 928 -468 936 -467
rect -481 -474 -473 -473
rect -405 -474 -397 -473
rect -330 -474 -322 -473
rect -253 -474 -245 -473
rect -176 -474 -168 -473
rect -100 -474 -92 -473
rect -9 -474 -1 -473
rect 71 -473 79 -472
rect 150 -472 158 -471
rect 226 -471 234 -470
rect 540 -470 548 -469
rect 622 -470 630 -469
rect 702 -470 710 -469
rect 1012 -470 1020 -469
rect 831 -471 839 -470
rect 928 -471 936 -470
rect 1012 -473 1020 -472
rect -481 -494 -473 -493
rect -405 -494 -397 -493
rect -330 -494 -322 -493
rect -253 -494 -245 -493
rect -176 -494 -168 -493
rect -100 -494 -92 -493
rect 540 -490 548 -489
rect 622 -490 630 -489
rect 702 -490 710 -489
rect 226 -491 234 -490
rect 150 -492 158 -491
rect 71 -493 79 -492
rect -9 -494 -1 -493
rect 831 -491 839 -490
rect 928 -491 936 -490
rect -481 -497 -473 -496
rect -405 -497 -397 -496
rect -330 -497 -322 -496
rect -253 -497 -245 -496
rect -176 -497 -168 -496
rect -100 -497 -92 -496
rect -9 -497 -1 -496
rect 71 -496 79 -495
rect 150 -495 158 -494
rect 226 -494 234 -493
rect 540 -493 548 -492
rect 622 -493 630 -492
rect 702 -493 710 -492
rect 1012 -493 1020 -492
rect 831 -494 839 -493
rect 928 -494 936 -493
rect 1012 -496 1020 -495
rect -481 -527 -473 -526
rect -405 -527 -397 -526
rect -330 -527 -322 -526
rect -253 -527 -245 -526
rect -176 -527 -168 -526
rect -100 -527 -92 -526
rect 540 -523 548 -522
rect 622 -523 630 -522
rect 702 -523 710 -522
rect 226 -524 234 -523
rect 150 -525 158 -524
rect 71 -526 79 -525
rect -9 -527 -1 -526
rect 831 -524 839 -523
rect 928 -524 936 -523
rect -481 -530 -473 -529
rect -405 -530 -397 -529
rect -330 -530 -322 -529
rect -253 -530 -245 -529
rect -176 -530 -168 -529
rect -100 -530 -92 -529
rect -9 -530 -1 -529
rect 71 -529 79 -528
rect 150 -528 158 -527
rect 226 -527 234 -526
rect 540 -526 548 -525
rect 622 -526 630 -525
rect 702 -526 710 -525
rect 1012 -526 1020 -525
rect 831 -527 839 -526
rect 928 -527 936 -526
rect 1012 -529 1020 -528
rect -481 -550 -473 -549
rect -405 -550 -397 -549
rect -330 -550 -322 -549
rect -253 -550 -245 -549
rect -176 -550 -168 -549
rect -100 -550 -92 -549
rect 540 -546 548 -545
rect 622 -546 630 -545
rect 702 -546 710 -545
rect 226 -547 234 -546
rect 150 -548 158 -547
rect 71 -549 79 -548
rect -9 -550 -1 -549
rect 831 -547 839 -546
rect 928 -547 936 -546
rect -481 -553 -473 -552
rect -405 -553 -397 -552
rect -330 -553 -322 -552
rect -253 -553 -245 -552
rect -176 -553 -168 -552
rect -100 -553 -92 -552
rect -9 -553 -1 -552
rect 71 -552 79 -551
rect 150 -551 158 -550
rect 226 -550 234 -549
rect 540 -549 548 -548
rect 622 -549 630 -548
rect 702 -549 710 -548
rect 1012 -549 1020 -548
rect 831 -550 839 -549
rect 928 -550 936 -549
rect 1012 -552 1020 -551
rect 869 -632 870 -624
rect 872 -632 873 -624
rect 892 -632 893 -624
rect 895 -632 896 -624
rect 466 -658 467 -650
rect 469 -658 470 -650
rect 489 -658 490 -650
rect 492 -658 493 -650
rect 64 -678 65 -670
rect 67 -678 68 -670
rect 87 -678 88 -670
rect 90 -678 91 -670
rect 943 -662 944 -654
rect 946 -662 947 -654
rect 966 -662 967 -654
rect 969 -662 970 -654
rect 540 -688 541 -680
rect 543 -688 544 -680
rect 563 -688 564 -680
rect 566 -688 567 -680
rect 677 -686 678 -678
rect 680 -686 681 -678
rect 700 -686 701 -678
rect 703 -686 704 -678
rect 734 -686 735 -678
rect 737 -686 738 -678
rect 757 -686 758 -678
rect 760 -686 761 -678
rect 814 -684 815 -676
rect 817 -684 818 -676
rect 837 -684 838 -676
rect 840 -684 841 -676
rect 138 -708 139 -700
rect 141 -708 142 -700
rect 161 -708 162 -700
rect 164 -708 165 -700
rect -371 -717 -363 -716
rect -371 -720 -363 -719
rect -128 -732 -127 -724
rect -125 -732 -124 -724
rect -105 -732 -104 -724
rect -102 -732 -101 -724
rect -71 -732 -70 -724
rect -68 -732 -67 -724
rect -48 -732 -47 -724
rect -45 -732 -44 -724
rect 9 -730 10 -722
rect 12 -730 13 -722
rect 32 -730 33 -722
rect 35 -730 36 -722
rect -371 -740 -363 -739
rect -460 -745 -452 -744
rect -371 -743 -363 -742
rect -460 -748 -452 -747
rect 274 -712 275 -704
rect 277 -712 278 -704
rect 297 -712 298 -704
rect 300 -712 301 -704
rect 331 -712 332 -704
rect 334 -712 335 -704
rect 354 -712 355 -704
rect 357 -712 358 -704
rect 411 -710 412 -702
rect 414 -710 415 -702
rect 434 -710 435 -702
rect 437 -710 438 -702
rect 877 -707 878 -699
rect 880 -707 881 -699
rect 900 -707 901 -699
rect 903 -707 904 -699
rect 474 -733 475 -725
rect 477 -733 478 -725
rect 497 -733 498 -725
rect 500 -733 501 -725
rect 72 -753 73 -745
rect 75 -753 76 -745
rect 95 -753 96 -745
rect 98 -753 99 -745
rect -460 -768 -452 -767
rect -460 -771 -452 -770
rect -319 -772 -311 -771
rect -319 -775 -311 -774
rect -394 -780 -386 -779
rect -394 -783 -386 -782
rect -319 -795 -311 -794
rect -460 -802 -452 -801
rect -319 -798 -311 -797
rect -394 -803 -386 -802
rect -460 -805 -452 -804
rect -394 -806 -386 -805
rect -460 -825 -452 -824
rect -460 -828 -452 -827
rect -349 -846 -341 -845
rect -349 -849 -341 -848
rect -349 -869 -341 -868
rect -349 -872 -341 -871
rect -521 -928 -513 -927
rect -455 -928 -447 -927
rect -63 -928 -55 -927
rect -366 -929 -358 -928
rect -521 -931 -513 -930
rect -455 -931 -447 -930
rect -366 -932 -358 -931
rect -63 -931 -55 -930
rect -521 -951 -513 -950
rect -455 -951 -447 -950
rect 270 -947 278 -946
rect -63 -951 -55 -950
rect -366 -952 -358 -951
rect -521 -954 -513 -953
rect -455 -954 -447 -953
rect -366 -955 -358 -954
rect -152 -956 -144 -955
rect -63 -954 -55 -953
rect 270 -950 278 -949
rect -152 -959 -144 -958
rect 270 -970 278 -969
rect 181 -975 189 -974
rect 270 -973 278 -972
rect -152 -979 -144 -978
rect -314 -984 -306 -983
rect -455 -985 -447 -984
rect -152 -982 -144 -981
rect 181 -978 189 -977
rect -11 -983 -3 -982
rect -455 -988 -447 -987
rect -314 -987 -306 -986
rect -11 -986 -3 -985
rect 813 -986 821 -985
rect -86 -991 -78 -990
rect -389 -992 -381 -991
rect 813 -989 821 -988
rect -389 -995 -381 -994
rect -86 -994 -78 -993
rect 181 -998 189 -997
rect 181 -1001 189 -1000
rect 322 -1002 330 -1001
rect -11 -1006 -3 -1005
rect -314 -1007 -306 -1006
rect -455 -1008 -447 -1007
rect -534 -1009 -526 -1008
rect -534 -1012 -526 -1011
rect -455 -1011 -447 -1010
rect -314 -1010 -306 -1009
rect -152 -1013 -144 -1012
rect -389 -1015 -381 -1014
rect -11 -1009 -3 -1008
rect 322 -1005 330 -1004
rect 813 -1009 821 -1008
rect 247 -1010 255 -1009
rect -86 -1014 -78 -1013
rect -389 -1018 -381 -1017
rect -152 -1016 -144 -1015
rect -86 -1017 -78 -1016
rect 247 -1013 255 -1012
rect 724 -1014 732 -1013
rect 813 -1012 821 -1011
rect 724 -1017 732 -1016
rect 322 -1025 330 -1024
rect -534 -1032 -526 -1031
rect -534 -1035 -526 -1034
rect 181 -1032 189 -1031
rect 322 -1028 330 -1027
rect 247 -1033 255 -1032
rect -152 -1036 -144 -1035
rect -152 -1039 -144 -1038
rect 181 -1035 189 -1034
rect 247 -1036 255 -1035
rect 724 -1037 732 -1036
rect 724 -1040 732 -1039
rect 865 -1041 873 -1040
rect 865 -1044 873 -1043
rect 790 -1049 798 -1048
rect -442 -1053 -434 -1052
rect -442 -1056 -434 -1055
rect 181 -1055 189 -1054
rect -41 -1057 -33 -1056
rect 790 -1052 798 -1051
rect -344 -1058 -336 -1057
rect -344 -1061 -336 -1060
rect -41 -1060 -33 -1059
rect 181 -1058 189 -1057
rect 865 -1064 873 -1063
rect 724 -1071 732 -1070
rect -442 -1076 -434 -1075
rect -442 -1079 -434 -1078
rect 865 -1067 873 -1066
rect 790 -1072 798 -1071
rect 292 -1076 300 -1075
rect 724 -1074 732 -1073
rect -41 -1080 -33 -1079
rect -344 -1081 -336 -1080
rect -344 -1084 -336 -1083
rect -41 -1083 -33 -1082
rect 292 -1079 300 -1078
rect 790 -1075 798 -1074
rect 724 -1094 732 -1093
rect 292 -1099 300 -1098
rect 724 -1097 732 -1096
rect 292 -1102 300 -1101
rect 835 -1115 843 -1114
rect 835 -1118 843 -1117
rect -213 -1139 -205 -1138
rect -147 -1139 -139 -1138
rect 835 -1138 843 -1137
rect -58 -1140 -50 -1139
rect -213 -1142 -205 -1141
rect -147 -1142 -139 -1141
rect -58 -1143 -50 -1142
rect 835 -1141 843 -1140
rect -213 -1162 -205 -1161
rect 120 -1158 128 -1157
rect 186 -1158 194 -1157
rect -147 -1162 -139 -1161
rect 275 -1159 283 -1158
rect -58 -1163 -50 -1162
rect -213 -1165 -205 -1164
rect -147 -1165 -139 -1164
rect 120 -1161 128 -1160
rect 186 -1161 194 -1160
rect -58 -1166 -50 -1165
rect 275 -1162 283 -1161
rect 120 -1181 128 -1180
rect 186 -1181 194 -1180
rect 275 -1182 283 -1181
rect 120 -1184 128 -1183
rect 186 -1184 194 -1183
rect 275 -1185 283 -1184
rect -6 -1195 2 -1194
rect -147 -1196 -139 -1195
rect 663 -1197 671 -1196
rect 729 -1197 737 -1196
rect -147 -1199 -139 -1198
rect -6 -1198 2 -1197
rect 818 -1198 826 -1197
rect -81 -1203 -73 -1202
rect 663 -1200 671 -1199
rect 729 -1200 737 -1199
rect 818 -1201 826 -1200
rect -81 -1206 -73 -1205
rect 327 -1214 335 -1213
rect 186 -1215 194 -1214
rect -6 -1218 2 -1217
rect -147 -1219 -139 -1218
rect -226 -1220 -218 -1219
rect -226 -1223 -218 -1222
rect -147 -1222 -139 -1221
rect -6 -1221 2 -1220
rect 186 -1218 194 -1217
rect 327 -1217 335 -1216
rect 663 -1220 671 -1219
rect 729 -1220 737 -1219
rect 252 -1222 260 -1221
rect 818 -1221 826 -1220
rect -81 -1226 -73 -1225
rect -81 -1229 -73 -1228
rect 252 -1225 260 -1224
rect 663 -1223 671 -1222
rect 729 -1223 737 -1222
rect 818 -1224 826 -1223
rect 327 -1237 335 -1236
rect 186 -1238 194 -1237
rect 107 -1239 115 -1238
rect -226 -1243 -218 -1242
rect -226 -1246 -218 -1245
rect 107 -1242 115 -1241
rect 186 -1241 194 -1240
rect 327 -1240 335 -1239
rect 252 -1245 260 -1244
rect 252 -1248 260 -1247
rect 870 -1253 878 -1252
rect 729 -1254 737 -1253
rect 729 -1257 737 -1256
rect 870 -1256 878 -1255
rect 795 -1261 803 -1260
rect 107 -1262 115 -1261
rect -134 -1264 -126 -1263
rect -134 -1267 -126 -1266
rect -36 -1269 -28 -1268
rect 107 -1265 115 -1264
rect 795 -1264 803 -1263
rect -36 -1272 -28 -1271
rect 870 -1276 878 -1275
rect 729 -1277 737 -1276
rect 650 -1278 658 -1277
rect 199 -1283 207 -1282
rect -134 -1287 -126 -1286
rect -134 -1290 -126 -1289
rect 199 -1286 207 -1285
rect 650 -1281 658 -1280
rect 729 -1280 737 -1279
rect 870 -1279 878 -1278
rect 795 -1284 803 -1283
rect 297 -1288 305 -1287
rect -36 -1292 -28 -1291
rect -36 -1295 -28 -1294
rect 297 -1291 305 -1290
rect 795 -1287 803 -1286
rect 650 -1301 658 -1300
rect 199 -1306 207 -1305
rect 199 -1309 207 -1308
rect 650 -1304 658 -1303
rect 297 -1311 305 -1310
rect 297 -1314 305 -1313
rect 742 -1322 750 -1321
rect 742 -1325 750 -1324
rect 840 -1327 848 -1326
rect 840 -1330 848 -1329
rect 742 -1345 750 -1344
rect 742 -1348 750 -1347
rect 840 -1350 848 -1349
rect 840 -1353 848 -1352
rect 516 -1509 524 -1508
rect 516 -1512 524 -1511
rect 516 -1532 524 -1531
rect 427 -1537 435 -1536
rect 516 -1535 524 -1534
rect 427 -1540 435 -1539
rect -127 -1557 -119 -1556
rect -127 -1560 -119 -1559
rect 427 -1560 435 -1559
rect 213 -1567 221 -1566
rect 427 -1563 435 -1562
rect 568 -1564 576 -1563
rect 213 -1570 221 -1569
rect 568 -1567 576 -1566
rect 493 -1572 501 -1571
rect 493 -1575 501 -1574
rect -127 -1580 -119 -1579
rect -216 -1585 -208 -1584
rect -127 -1583 -119 -1582
rect -216 -1588 -208 -1587
rect 568 -1587 576 -1586
rect 213 -1590 221 -1589
rect 124 -1595 132 -1594
rect 213 -1593 221 -1592
rect 427 -1594 435 -1593
rect 568 -1590 576 -1589
rect 493 -1595 501 -1594
rect 124 -1598 132 -1597
rect 427 -1597 435 -1596
rect 493 -1598 501 -1597
rect -216 -1608 -208 -1607
rect -432 -1613 -424 -1612
rect -216 -1611 -208 -1610
rect -75 -1612 -67 -1611
rect -432 -1616 -424 -1615
rect -75 -1615 -67 -1614
rect 427 -1617 435 -1616
rect 124 -1618 132 -1617
rect -150 -1620 -142 -1619
rect -150 -1623 -142 -1622
rect 124 -1621 132 -1620
rect 265 -1622 273 -1621
rect 427 -1620 435 -1619
rect 265 -1625 273 -1624
rect 190 -1630 198 -1629
rect -75 -1635 -67 -1634
rect -432 -1636 -424 -1635
rect 190 -1633 198 -1632
rect -521 -1641 -513 -1640
rect -432 -1639 -424 -1638
rect -216 -1642 -208 -1641
rect -521 -1644 -513 -1643
rect -75 -1638 -67 -1637
rect 538 -1638 546 -1637
rect -150 -1643 -142 -1642
rect -216 -1645 -208 -1644
rect 265 -1645 273 -1644
rect 538 -1641 546 -1640
rect -150 -1646 -142 -1645
rect 124 -1652 132 -1651
rect 265 -1648 273 -1647
rect 190 -1653 198 -1652
rect 124 -1655 132 -1654
rect 190 -1656 198 -1655
rect -521 -1664 -513 -1663
rect -521 -1667 -513 -1666
rect 538 -1661 546 -1660
rect -216 -1665 -208 -1664
rect -380 -1668 -372 -1667
rect -380 -1671 -372 -1670
rect -216 -1668 -208 -1667
rect 538 -1664 546 -1663
rect 124 -1675 132 -1674
rect -455 -1676 -447 -1675
rect -455 -1679 -447 -1678
rect 124 -1678 132 -1677
rect -105 -1686 -97 -1685
rect -380 -1691 -372 -1690
rect -105 -1689 -97 -1688
rect -521 -1698 -513 -1697
rect -380 -1694 -372 -1693
rect 235 -1696 243 -1695
rect -455 -1699 -447 -1698
rect -521 -1701 -513 -1700
rect -455 -1702 -447 -1701
rect 235 -1699 243 -1698
rect -105 -1709 -97 -1708
rect -105 -1712 -97 -1711
rect 235 -1719 243 -1718
rect -521 -1721 -513 -1720
rect 366 -1720 374 -1719
rect 432 -1720 440 -1719
rect -521 -1724 -513 -1723
rect 235 -1722 243 -1721
rect 521 -1721 529 -1720
rect 366 -1723 374 -1722
rect 432 -1723 440 -1722
rect 521 -1724 529 -1723
rect -410 -1742 -402 -1741
rect 366 -1743 374 -1742
rect 432 -1743 440 -1742
rect -410 -1745 -402 -1744
rect 521 -1744 529 -1743
rect 366 -1746 374 -1745
rect 432 -1746 440 -1745
rect 521 -1747 529 -1746
rect -410 -1765 -402 -1764
rect -410 -1768 -402 -1767
rect -277 -1768 -269 -1767
rect -211 -1768 -203 -1767
rect -122 -1769 -114 -1768
rect -277 -1771 -269 -1770
rect -211 -1771 -203 -1770
rect -122 -1772 -114 -1771
rect 63 -1778 71 -1777
rect 129 -1778 137 -1777
rect 573 -1776 581 -1775
rect 432 -1777 440 -1776
rect 218 -1779 226 -1778
rect 63 -1781 71 -1780
rect 129 -1781 137 -1780
rect 218 -1782 226 -1781
rect 432 -1780 440 -1779
rect 573 -1779 581 -1778
rect 498 -1784 506 -1783
rect -277 -1791 -269 -1790
rect -211 -1791 -203 -1790
rect 498 -1787 506 -1786
rect -122 -1792 -114 -1791
rect -277 -1794 -269 -1793
rect -211 -1794 -203 -1793
rect -122 -1795 -114 -1794
rect 63 -1801 71 -1800
rect 129 -1801 137 -1800
rect 573 -1799 581 -1798
rect 432 -1800 440 -1799
rect 353 -1801 361 -1800
rect 218 -1802 226 -1801
rect 63 -1804 71 -1803
rect 129 -1804 137 -1803
rect 218 -1805 226 -1804
rect 353 -1804 361 -1803
rect 432 -1803 440 -1802
rect 573 -1802 581 -1801
rect 498 -1807 506 -1806
rect 498 -1810 506 -1809
rect -582 -1824 -574 -1823
rect -516 -1824 -508 -1823
rect -427 -1825 -419 -1824
rect -70 -1824 -62 -1823
rect 353 -1824 361 -1823
rect -211 -1825 -203 -1824
rect -582 -1827 -574 -1826
rect -516 -1827 -508 -1826
rect -427 -1828 -419 -1827
rect -211 -1828 -203 -1827
rect -70 -1827 -62 -1826
rect -145 -1832 -137 -1831
rect -145 -1835 -137 -1834
rect 353 -1827 361 -1826
rect 270 -1834 278 -1833
rect 129 -1835 137 -1834
rect 129 -1838 137 -1837
rect 270 -1837 278 -1836
rect 195 -1842 203 -1841
rect -582 -1847 -574 -1846
rect -516 -1847 -508 -1846
rect -427 -1848 -419 -1847
rect -582 -1850 -574 -1849
rect -516 -1850 -508 -1849
rect -70 -1847 -62 -1846
rect -211 -1848 -203 -1847
rect -290 -1849 -282 -1848
rect -427 -1851 -419 -1850
rect 195 -1845 203 -1844
rect 445 -1845 453 -1844
rect -290 -1852 -282 -1851
rect -211 -1851 -203 -1850
rect -70 -1850 -62 -1849
rect 445 -1848 453 -1847
rect 543 -1850 551 -1849
rect -145 -1855 -137 -1854
rect -145 -1858 -137 -1857
rect 270 -1857 278 -1856
rect 543 -1853 551 -1852
rect 129 -1858 137 -1857
rect 50 -1859 58 -1858
rect 50 -1862 58 -1861
rect 129 -1861 137 -1860
rect 270 -1860 278 -1859
rect 195 -1865 203 -1864
rect -290 -1872 -282 -1871
rect 195 -1868 203 -1867
rect 445 -1868 453 -1867
rect -290 -1875 -282 -1874
rect 445 -1871 453 -1870
rect 543 -1873 551 -1872
rect -375 -1880 -367 -1879
rect -516 -1881 -508 -1880
rect 543 -1876 551 -1875
rect 50 -1882 58 -1881
rect -516 -1884 -508 -1883
rect -375 -1883 -367 -1882
rect -450 -1888 -442 -1887
rect -450 -1891 -442 -1890
rect 50 -1885 58 -1884
rect -198 -1893 -190 -1892
rect -198 -1896 -190 -1895
rect -100 -1898 -92 -1897
rect -375 -1903 -367 -1902
rect -516 -1904 -508 -1903
rect -595 -1905 -587 -1904
rect -100 -1901 -92 -1900
rect 142 -1903 150 -1902
rect -595 -1908 -587 -1907
rect -516 -1907 -508 -1906
rect -375 -1906 -367 -1905
rect 142 -1906 150 -1905
rect 240 -1908 248 -1907
rect -450 -1911 -442 -1910
rect -450 -1914 -442 -1913
rect 240 -1911 248 -1910
rect -198 -1916 -190 -1915
rect -198 -1919 -190 -1918
rect -100 -1921 -92 -1920
rect -595 -1928 -587 -1927
rect -100 -1924 -92 -1923
rect 142 -1926 150 -1925
rect -595 -1931 -587 -1930
rect 142 -1929 150 -1928
rect 240 -1931 248 -1930
rect 240 -1934 248 -1933
rect -503 -1949 -495 -1948
rect -503 -1952 -495 -1951
rect -405 -1954 -397 -1953
rect -405 -1957 -397 -1956
rect -503 -1972 -495 -1971
rect -503 -1975 -495 -1974
rect -405 -1977 -397 -1976
rect -405 -1980 -397 -1979
rect 450 -2047 451 -2039
rect 453 -2047 454 -2039
rect 473 -2047 474 -2039
rect 476 -2047 477 -2039
rect 524 -2077 525 -2069
rect 527 -2077 528 -2069
rect 547 -2077 548 -2069
rect 550 -2077 551 -2069
rect 258 -2101 259 -2093
rect 261 -2101 262 -2093
rect 281 -2101 282 -2093
rect 284 -2101 285 -2093
rect 315 -2101 316 -2093
rect 318 -2101 319 -2093
rect 338 -2101 339 -2093
rect 341 -2101 342 -2093
rect 395 -2099 396 -2091
rect 398 -2099 399 -2091
rect 418 -2099 419 -2091
rect 421 -2099 422 -2091
rect 458 -2122 459 -2114
rect 461 -2122 462 -2114
rect 481 -2122 482 -2114
rect 484 -2122 485 -2114
<< ndcontact >>
rect -513 -470 -507 -466
rect -437 -470 -431 -466
rect -362 -470 -356 -466
rect -285 -470 -279 -466
rect -208 -470 -202 -466
rect -132 -470 -126 -466
rect -41 -470 -35 -466
rect 39 -469 45 -465
rect 118 -468 124 -464
rect 194 -467 200 -463
rect 508 -466 514 -462
rect 590 -466 596 -462
rect 670 -466 676 -462
rect 799 -467 805 -463
rect 896 -467 902 -463
rect -513 -478 -507 -474
rect -437 -478 -431 -474
rect -362 -478 -356 -474
rect -285 -478 -279 -474
rect -208 -478 -202 -474
rect -132 -478 -126 -474
rect -41 -478 -35 -474
rect 39 -477 45 -473
rect 118 -476 124 -472
rect 194 -475 200 -471
rect 508 -474 514 -470
rect 590 -474 596 -470
rect 670 -474 676 -470
rect 980 -469 986 -465
rect 799 -475 805 -471
rect 896 -475 902 -471
rect 980 -477 986 -473
rect -513 -493 -507 -489
rect -437 -493 -431 -489
rect -362 -493 -356 -489
rect -285 -493 -279 -489
rect -208 -493 -202 -489
rect -132 -493 -126 -489
rect -41 -493 -35 -489
rect 39 -492 45 -488
rect 118 -491 124 -487
rect 194 -490 200 -486
rect 508 -489 514 -485
rect 590 -489 596 -485
rect 670 -489 676 -485
rect 799 -490 805 -486
rect 896 -490 902 -486
rect -513 -501 -507 -497
rect -437 -501 -431 -497
rect -362 -501 -356 -497
rect -285 -501 -279 -497
rect -208 -501 -202 -497
rect -132 -501 -126 -497
rect -41 -501 -35 -497
rect 39 -500 45 -496
rect 118 -499 124 -495
rect 194 -498 200 -494
rect 508 -497 514 -493
rect 590 -497 596 -493
rect 670 -497 676 -493
rect 980 -492 986 -488
rect 799 -498 805 -494
rect 896 -498 902 -494
rect 980 -500 986 -496
rect -513 -526 -507 -522
rect -437 -526 -431 -522
rect -362 -526 -356 -522
rect -285 -526 -279 -522
rect -208 -526 -202 -522
rect -132 -526 -126 -522
rect -41 -526 -35 -522
rect 39 -525 45 -521
rect 118 -524 124 -520
rect 194 -523 200 -519
rect 508 -522 514 -518
rect 590 -522 596 -518
rect 670 -522 676 -518
rect 799 -523 805 -519
rect 896 -523 902 -519
rect -513 -534 -507 -530
rect -437 -534 -431 -530
rect -362 -534 -356 -530
rect -285 -534 -279 -530
rect -208 -534 -202 -530
rect -132 -534 -126 -530
rect -41 -534 -35 -530
rect 39 -533 45 -529
rect 118 -532 124 -528
rect 194 -531 200 -527
rect 508 -530 514 -526
rect 590 -530 596 -526
rect 670 -530 676 -526
rect 980 -525 986 -521
rect 799 -531 805 -527
rect 896 -531 902 -527
rect 980 -533 986 -529
rect -513 -549 -507 -545
rect -437 -549 -431 -545
rect -362 -549 -356 -545
rect -285 -549 -279 -545
rect -208 -549 -202 -545
rect -132 -549 -126 -545
rect -41 -549 -35 -545
rect 39 -548 45 -544
rect 118 -547 124 -543
rect 194 -546 200 -542
rect 508 -545 514 -541
rect 590 -545 596 -541
rect 670 -545 676 -541
rect 799 -546 805 -542
rect 896 -546 902 -542
rect -513 -557 -507 -553
rect -437 -557 -431 -553
rect -362 -557 -356 -553
rect -285 -557 -279 -553
rect -208 -557 -202 -553
rect -132 -557 -126 -553
rect -41 -557 -35 -553
rect 39 -556 45 -552
rect 118 -555 124 -551
rect 194 -554 200 -550
rect 508 -553 514 -549
rect 590 -553 596 -549
rect 670 -553 676 -549
rect 980 -548 986 -544
rect 799 -554 805 -550
rect 896 -554 902 -550
rect 980 -556 986 -552
rect 865 -664 869 -658
rect 873 -664 877 -658
rect 888 -664 892 -658
rect 896 -664 900 -658
rect 462 -690 466 -684
rect 470 -690 474 -684
rect 485 -690 489 -684
rect 493 -690 497 -684
rect 60 -710 64 -704
rect 68 -710 72 -704
rect 83 -710 87 -704
rect 91 -710 95 -704
rect -403 -716 -397 -712
rect -403 -724 -397 -720
rect -403 -739 -397 -735
rect -492 -744 -486 -740
rect -403 -747 -397 -743
rect -492 -752 -486 -748
rect 134 -740 138 -734
rect 142 -740 146 -734
rect 157 -740 161 -734
rect 165 -740 169 -734
rect 939 -694 943 -688
rect 947 -694 951 -688
rect 962 -694 966 -688
rect 970 -694 974 -688
rect 536 -720 540 -714
rect 544 -720 548 -714
rect 559 -720 563 -714
rect 567 -720 571 -714
rect 673 -718 677 -712
rect 681 -718 685 -712
rect 696 -718 700 -712
rect 704 -718 708 -712
rect 730 -718 734 -712
rect 738 -718 742 -712
rect 753 -718 757 -712
rect 761 -718 765 -712
rect 810 -716 814 -710
rect 818 -716 822 -710
rect 833 -716 837 -710
rect 841 -716 845 -710
rect 270 -744 274 -738
rect 278 -744 282 -738
rect 293 -744 297 -738
rect 301 -744 305 -738
rect 327 -744 331 -738
rect 335 -744 339 -738
rect 350 -744 354 -738
rect 358 -744 362 -738
rect 407 -742 411 -736
rect 415 -742 419 -736
rect 430 -742 434 -736
rect 438 -742 442 -736
rect -492 -767 -486 -763
rect -132 -764 -128 -758
rect -124 -764 -120 -758
rect -109 -764 -105 -758
rect -101 -764 -97 -758
rect -75 -764 -71 -758
rect -67 -764 -63 -758
rect -52 -764 -48 -758
rect -44 -764 -40 -758
rect 5 -762 9 -756
rect 13 -762 17 -756
rect 28 -762 32 -756
rect 36 -762 40 -756
rect -492 -775 -486 -771
rect -351 -771 -345 -767
rect -426 -779 -420 -775
rect -351 -779 -345 -775
rect 873 -739 877 -733
rect 881 -739 885 -733
rect 896 -739 900 -733
rect 904 -739 908 -733
rect 470 -765 474 -759
rect 478 -765 482 -759
rect 493 -765 497 -759
rect 501 -765 505 -759
rect -426 -787 -420 -783
rect 68 -785 72 -779
rect 76 -785 80 -779
rect 91 -785 95 -779
rect 99 -785 103 -779
rect -351 -794 -345 -790
rect -492 -801 -486 -797
rect -426 -802 -420 -798
rect -351 -802 -345 -798
rect -492 -809 -486 -805
rect -426 -810 -420 -806
rect -492 -824 -486 -820
rect -492 -832 -486 -828
rect -381 -845 -375 -841
rect -381 -853 -375 -849
rect -381 -868 -375 -864
rect -381 -876 -375 -872
rect -553 -927 -547 -923
rect -487 -927 -481 -923
rect -398 -928 -392 -924
rect -95 -927 -89 -923
rect -553 -935 -547 -931
rect -487 -935 -481 -931
rect -398 -936 -392 -932
rect -95 -935 -89 -931
rect 238 -946 244 -942
rect -553 -950 -547 -946
rect -487 -950 -481 -946
rect -398 -951 -392 -947
rect -95 -950 -89 -946
rect -553 -958 -547 -954
rect -487 -958 -481 -954
rect -398 -959 -392 -955
rect -184 -955 -178 -951
rect -95 -958 -89 -954
rect 238 -954 244 -950
rect -184 -963 -178 -959
rect 238 -969 244 -965
rect 149 -974 155 -970
rect -184 -978 -178 -974
rect 238 -977 244 -973
rect -487 -984 -481 -980
rect -346 -983 -340 -979
rect -184 -986 -178 -982
rect -43 -982 -37 -978
rect 149 -982 155 -978
rect 781 -985 787 -981
rect -487 -992 -481 -988
rect -421 -991 -415 -987
rect -346 -991 -340 -987
rect -118 -990 -112 -986
rect -43 -990 -37 -986
rect 781 -993 787 -989
rect -421 -999 -415 -995
rect -118 -998 -112 -994
rect 149 -997 155 -993
rect -566 -1008 -560 -1004
rect -487 -1007 -481 -1003
rect -346 -1006 -340 -1002
rect -43 -1005 -37 -1001
rect 149 -1005 155 -1001
rect 290 -1001 296 -997
rect -566 -1016 -560 -1012
rect -487 -1015 -481 -1011
rect -421 -1014 -415 -1010
rect -346 -1014 -340 -1010
rect -184 -1012 -178 -1008
rect -118 -1013 -112 -1009
rect -43 -1013 -37 -1009
rect 215 -1009 221 -1005
rect 290 -1009 296 -1005
rect 781 -1008 787 -1004
rect -421 -1022 -415 -1018
rect -184 -1020 -178 -1016
rect -118 -1021 -112 -1017
rect 215 -1017 221 -1013
rect 692 -1013 698 -1009
rect 781 -1016 787 -1012
rect 290 -1024 296 -1020
rect 692 -1021 698 -1017
rect -566 -1031 -560 -1027
rect 149 -1031 155 -1027
rect -566 -1039 -560 -1035
rect -184 -1035 -178 -1031
rect 215 -1032 221 -1028
rect 290 -1032 296 -1028
rect -184 -1043 -178 -1039
rect 149 -1039 155 -1035
rect 215 -1040 221 -1036
rect 692 -1036 698 -1032
rect 692 -1044 698 -1040
rect 833 -1040 839 -1036
rect 758 -1048 764 -1044
rect -474 -1052 -468 -1048
rect 833 -1048 839 -1044
rect -474 -1060 -468 -1056
rect -376 -1057 -370 -1053
rect -73 -1056 -67 -1052
rect 149 -1054 155 -1050
rect 758 -1056 764 -1052
rect -376 -1065 -370 -1061
rect -73 -1064 -67 -1060
rect 149 -1062 155 -1058
rect 833 -1063 839 -1059
rect 692 -1070 698 -1066
rect 758 -1071 764 -1067
rect -474 -1075 -468 -1071
rect 260 -1075 266 -1071
rect -474 -1083 -468 -1079
rect -376 -1080 -370 -1076
rect -73 -1079 -67 -1075
rect 833 -1071 839 -1067
rect 692 -1078 698 -1074
rect -376 -1088 -370 -1084
rect -73 -1087 -67 -1083
rect 260 -1083 266 -1079
rect 758 -1079 764 -1075
rect 692 -1093 698 -1089
rect 260 -1098 266 -1094
rect 692 -1101 698 -1097
rect 260 -1106 266 -1102
rect 803 -1114 809 -1110
rect 803 -1122 809 -1118
rect -245 -1138 -239 -1134
rect -179 -1138 -173 -1134
rect -90 -1139 -84 -1135
rect 803 -1137 809 -1133
rect -245 -1146 -239 -1142
rect -179 -1146 -173 -1142
rect -90 -1147 -84 -1143
rect 803 -1145 809 -1141
rect 88 -1157 94 -1153
rect -245 -1161 -239 -1157
rect -179 -1161 -173 -1157
rect 154 -1157 160 -1153
rect 243 -1158 249 -1154
rect -90 -1162 -84 -1158
rect -245 -1169 -239 -1165
rect -179 -1169 -173 -1165
rect 88 -1165 94 -1161
rect 154 -1165 160 -1161
rect -90 -1170 -84 -1166
rect 243 -1166 249 -1162
rect 88 -1180 94 -1176
rect 154 -1180 160 -1176
rect 243 -1181 249 -1177
rect 88 -1188 94 -1184
rect 154 -1188 160 -1184
rect 243 -1189 249 -1185
rect -179 -1195 -173 -1191
rect -38 -1194 -32 -1190
rect 631 -1196 637 -1192
rect 697 -1196 703 -1192
rect 786 -1197 792 -1193
rect -179 -1203 -173 -1199
rect -113 -1202 -107 -1198
rect -38 -1202 -32 -1198
rect 631 -1204 637 -1200
rect 697 -1204 703 -1200
rect 786 -1205 792 -1201
rect -113 -1210 -107 -1206
rect -258 -1219 -252 -1215
rect -179 -1218 -173 -1214
rect -38 -1217 -32 -1213
rect 154 -1214 160 -1210
rect 295 -1213 301 -1209
rect -258 -1227 -252 -1223
rect -179 -1226 -173 -1222
rect -113 -1225 -107 -1221
rect -38 -1225 -32 -1221
rect 154 -1222 160 -1218
rect 220 -1221 226 -1217
rect 295 -1221 301 -1217
rect 631 -1219 637 -1215
rect 697 -1219 703 -1215
rect 786 -1220 792 -1216
rect -113 -1233 -107 -1229
rect 220 -1229 226 -1225
rect 631 -1227 637 -1223
rect 697 -1227 703 -1223
rect 786 -1228 792 -1224
rect 75 -1238 81 -1234
rect -258 -1242 -252 -1238
rect 154 -1237 160 -1233
rect 295 -1236 301 -1232
rect -258 -1250 -252 -1246
rect 75 -1246 81 -1242
rect 154 -1245 160 -1241
rect 220 -1244 226 -1240
rect 295 -1244 301 -1240
rect 220 -1252 226 -1248
rect 697 -1253 703 -1249
rect 838 -1252 844 -1248
rect -166 -1263 -160 -1259
rect 75 -1261 81 -1257
rect 697 -1261 703 -1257
rect 763 -1260 769 -1256
rect 838 -1260 844 -1256
rect -166 -1271 -160 -1267
rect -68 -1268 -62 -1264
rect 75 -1269 81 -1265
rect 763 -1268 769 -1264
rect -68 -1276 -62 -1272
rect 618 -1277 624 -1273
rect 697 -1276 703 -1272
rect 838 -1275 844 -1271
rect 167 -1282 173 -1278
rect -166 -1286 -160 -1282
rect -166 -1294 -160 -1290
rect -68 -1291 -62 -1287
rect 167 -1290 173 -1286
rect 265 -1287 271 -1283
rect 618 -1285 624 -1281
rect 697 -1284 703 -1280
rect 763 -1283 769 -1279
rect 838 -1283 844 -1279
rect -68 -1299 -62 -1295
rect 265 -1295 271 -1291
rect 763 -1291 769 -1287
rect 618 -1300 624 -1296
rect 167 -1305 173 -1301
rect 167 -1313 173 -1309
rect 265 -1310 271 -1306
rect 618 -1308 624 -1304
rect 265 -1318 271 -1314
rect 710 -1321 716 -1317
rect 710 -1329 716 -1325
rect 808 -1326 814 -1322
rect 808 -1334 814 -1330
rect 710 -1344 716 -1340
rect 710 -1352 716 -1348
rect 808 -1349 814 -1345
rect 808 -1357 814 -1353
rect 484 -1508 490 -1504
rect 484 -1516 490 -1512
rect 484 -1531 490 -1527
rect 395 -1536 401 -1532
rect 484 -1539 490 -1535
rect 395 -1544 401 -1540
rect -159 -1556 -153 -1552
rect 395 -1559 401 -1555
rect -159 -1564 -153 -1560
rect 181 -1566 187 -1562
rect 395 -1567 401 -1563
rect 536 -1563 542 -1559
rect 181 -1574 187 -1570
rect 461 -1571 467 -1567
rect 536 -1571 542 -1567
rect -159 -1579 -153 -1575
rect 461 -1579 467 -1575
rect -248 -1584 -242 -1580
rect -159 -1587 -153 -1583
rect -248 -1592 -242 -1588
rect 181 -1589 187 -1585
rect 536 -1586 542 -1582
rect 92 -1594 98 -1590
rect 181 -1597 187 -1593
rect 395 -1593 401 -1589
rect 461 -1594 467 -1590
rect 536 -1594 542 -1590
rect 92 -1602 98 -1598
rect 395 -1601 401 -1597
rect 461 -1602 467 -1598
rect -248 -1607 -242 -1603
rect -464 -1612 -458 -1608
rect -248 -1615 -242 -1611
rect -107 -1611 -101 -1607
rect -464 -1620 -458 -1616
rect -182 -1619 -176 -1615
rect -107 -1619 -101 -1615
rect 92 -1617 98 -1613
rect 395 -1616 401 -1612
rect -182 -1627 -176 -1623
rect 92 -1625 98 -1621
rect 233 -1621 239 -1617
rect 395 -1624 401 -1620
rect 158 -1629 164 -1625
rect 233 -1629 239 -1625
rect -464 -1635 -458 -1631
rect -107 -1634 -101 -1630
rect -553 -1640 -547 -1636
rect 158 -1637 164 -1633
rect 506 -1637 512 -1633
rect -464 -1643 -458 -1639
rect -248 -1641 -242 -1637
rect -182 -1642 -176 -1638
rect -553 -1648 -547 -1644
rect -107 -1642 -101 -1638
rect -248 -1649 -242 -1645
rect 233 -1644 239 -1640
rect 506 -1645 512 -1641
rect -182 -1650 -176 -1646
rect 92 -1651 98 -1647
rect 158 -1652 164 -1648
rect 233 -1652 239 -1648
rect 92 -1659 98 -1655
rect -553 -1663 -547 -1659
rect 158 -1660 164 -1656
rect 506 -1660 512 -1656
rect -553 -1671 -547 -1667
rect -412 -1667 -406 -1663
rect -248 -1664 -242 -1660
rect -487 -1675 -481 -1671
rect -412 -1675 -406 -1671
rect -248 -1672 -242 -1668
rect 506 -1668 512 -1664
rect 92 -1674 98 -1670
rect -487 -1683 -481 -1679
rect -137 -1685 -131 -1681
rect 92 -1682 98 -1678
rect -412 -1690 -406 -1686
rect -137 -1693 -131 -1689
rect -553 -1697 -547 -1693
rect -487 -1698 -481 -1694
rect -412 -1698 -406 -1694
rect 203 -1695 209 -1691
rect -553 -1705 -547 -1701
rect -487 -1706 -481 -1702
rect 203 -1703 209 -1699
rect -137 -1708 -131 -1704
rect -137 -1716 -131 -1712
rect -553 -1720 -547 -1716
rect 203 -1718 209 -1714
rect 334 -1719 340 -1715
rect 400 -1719 406 -1715
rect 489 -1720 495 -1716
rect -553 -1728 -547 -1724
rect 203 -1726 209 -1722
rect 334 -1727 340 -1723
rect 400 -1727 406 -1723
rect 489 -1728 495 -1724
rect -442 -1741 -436 -1737
rect 334 -1742 340 -1738
rect 400 -1742 406 -1738
rect 489 -1743 495 -1739
rect -442 -1749 -436 -1745
rect 334 -1750 340 -1746
rect 400 -1750 406 -1746
rect 489 -1751 495 -1747
rect -442 -1764 -436 -1760
rect -309 -1767 -303 -1763
rect -442 -1772 -436 -1768
rect -243 -1767 -237 -1763
rect -154 -1768 -148 -1764
rect -309 -1775 -303 -1771
rect -243 -1775 -237 -1771
rect -154 -1776 -148 -1772
rect 31 -1777 37 -1773
rect 97 -1777 103 -1773
rect 186 -1778 192 -1774
rect 400 -1776 406 -1772
rect 541 -1775 547 -1771
rect 31 -1785 37 -1781
rect 97 -1785 103 -1781
rect 186 -1786 192 -1782
rect 400 -1784 406 -1780
rect 466 -1783 472 -1779
rect 541 -1783 547 -1779
rect -309 -1790 -303 -1786
rect -243 -1790 -237 -1786
rect -154 -1791 -148 -1787
rect 466 -1791 472 -1787
rect -309 -1798 -303 -1794
rect -243 -1798 -237 -1794
rect -154 -1799 -148 -1795
rect 31 -1800 37 -1796
rect 97 -1800 103 -1796
rect 186 -1801 192 -1797
rect 321 -1800 327 -1796
rect 400 -1799 406 -1795
rect 541 -1798 547 -1794
rect 31 -1808 37 -1804
rect 97 -1808 103 -1804
rect 186 -1809 192 -1805
rect 321 -1808 327 -1804
rect 400 -1807 406 -1803
rect 466 -1806 472 -1802
rect 541 -1806 547 -1802
rect 466 -1814 472 -1810
rect -614 -1823 -608 -1819
rect -548 -1823 -542 -1819
rect -459 -1824 -453 -1820
rect -243 -1824 -237 -1820
rect -102 -1823 -96 -1819
rect 321 -1823 327 -1819
rect -614 -1831 -608 -1827
rect -548 -1831 -542 -1827
rect -459 -1832 -453 -1828
rect -243 -1832 -237 -1828
rect -177 -1831 -171 -1827
rect -102 -1831 -96 -1827
rect 97 -1834 103 -1830
rect -177 -1839 -171 -1835
rect 238 -1833 244 -1829
rect 321 -1831 327 -1827
rect 97 -1842 103 -1838
rect 163 -1841 169 -1837
rect 238 -1841 244 -1837
rect -614 -1846 -608 -1842
rect -548 -1846 -542 -1842
rect -459 -1847 -453 -1843
rect -322 -1848 -316 -1844
rect -614 -1854 -608 -1850
rect -548 -1854 -542 -1850
rect -243 -1847 -237 -1843
rect -102 -1846 -96 -1842
rect 413 -1844 419 -1840
rect -459 -1855 -453 -1851
rect 163 -1849 169 -1845
rect -322 -1856 -316 -1852
rect -243 -1855 -237 -1851
rect -177 -1854 -171 -1850
rect -102 -1854 -96 -1850
rect 413 -1852 419 -1848
rect 511 -1849 517 -1845
rect -177 -1862 -171 -1858
rect 18 -1858 24 -1854
rect 97 -1857 103 -1853
rect 238 -1856 244 -1852
rect 511 -1857 517 -1853
rect 18 -1866 24 -1862
rect 97 -1865 103 -1861
rect 163 -1864 169 -1860
rect 238 -1864 244 -1860
rect 413 -1867 419 -1863
rect -322 -1871 -316 -1867
rect 163 -1872 169 -1868
rect -548 -1880 -542 -1876
rect -407 -1879 -401 -1875
rect -322 -1879 -316 -1875
rect 413 -1875 419 -1871
rect 511 -1872 517 -1868
rect 18 -1881 24 -1877
rect 511 -1880 517 -1876
rect -548 -1888 -542 -1884
rect -482 -1887 -476 -1883
rect -407 -1887 -401 -1883
rect -482 -1895 -476 -1891
rect -230 -1892 -224 -1888
rect 18 -1889 24 -1885
rect -627 -1904 -621 -1900
rect -548 -1903 -542 -1899
rect -407 -1902 -401 -1898
rect -230 -1900 -224 -1896
rect -132 -1897 -126 -1893
rect -132 -1905 -126 -1901
rect 110 -1902 116 -1898
rect -627 -1912 -621 -1908
rect -548 -1911 -542 -1907
rect -482 -1910 -476 -1906
rect -407 -1910 -401 -1906
rect 110 -1910 116 -1906
rect 208 -1907 214 -1903
rect -482 -1918 -476 -1914
rect -230 -1915 -224 -1911
rect 208 -1915 214 -1911
rect -230 -1923 -224 -1919
rect -132 -1920 -126 -1916
rect -627 -1927 -621 -1923
rect -132 -1928 -126 -1924
rect 110 -1925 116 -1921
rect -627 -1935 -621 -1931
rect 110 -1933 116 -1929
rect 208 -1930 214 -1926
rect 208 -1938 214 -1934
rect -535 -1948 -529 -1944
rect -535 -1956 -529 -1952
rect -437 -1953 -431 -1949
rect -437 -1961 -431 -1957
rect -535 -1971 -529 -1967
rect -535 -1979 -529 -1975
rect -437 -1976 -431 -1972
rect -437 -1984 -431 -1980
rect 446 -2079 450 -2073
rect 454 -2079 458 -2073
rect 469 -2079 473 -2073
rect 477 -2079 481 -2073
rect 520 -2109 524 -2103
rect 528 -2109 532 -2103
rect 543 -2109 547 -2103
rect 551 -2109 555 -2103
rect 254 -2133 258 -2127
rect 262 -2133 266 -2127
rect 277 -2133 281 -2127
rect 285 -2133 289 -2127
rect 311 -2133 315 -2127
rect 319 -2133 323 -2127
rect 334 -2133 338 -2127
rect 342 -2133 346 -2127
rect 391 -2131 395 -2125
rect 399 -2131 403 -2125
rect 414 -2131 418 -2125
rect 422 -2131 426 -2125
rect 454 -2154 458 -2148
rect 462 -2154 466 -2148
rect 477 -2154 481 -2148
rect 485 -2154 489 -2148
<< pdcontact >>
rect -481 -470 -473 -466
rect -405 -470 -397 -466
rect -330 -470 -322 -466
rect -253 -470 -245 -466
rect -176 -470 -168 -466
rect -100 -470 -92 -466
rect -9 -470 -1 -466
rect 71 -469 79 -465
rect 150 -468 158 -464
rect 226 -467 234 -463
rect 540 -466 548 -462
rect 622 -466 630 -462
rect 702 -466 710 -462
rect 831 -467 839 -463
rect 928 -467 936 -463
rect -481 -478 -473 -474
rect -405 -478 -397 -474
rect -330 -478 -322 -474
rect -253 -478 -245 -474
rect -176 -478 -168 -474
rect -100 -478 -92 -474
rect -9 -478 -1 -474
rect 71 -477 79 -473
rect 150 -476 158 -472
rect 226 -475 234 -471
rect 540 -474 548 -470
rect 622 -474 630 -470
rect 1012 -469 1020 -465
rect 702 -474 710 -470
rect 831 -475 839 -471
rect 928 -475 936 -471
rect 1012 -477 1020 -473
rect -481 -493 -473 -489
rect -405 -493 -397 -489
rect -330 -493 -322 -489
rect -253 -493 -245 -489
rect -176 -493 -168 -489
rect -100 -493 -92 -489
rect -9 -493 -1 -489
rect 71 -492 79 -488
rect 150 -491 158 -487
rect 226 -490 234 -486
rect 540 -489 548 -485
rect 622 -489 630 -485
rect 702 -489 710 -485
rect 831 -490 839 -486
rect 928 -490 936 -486
rect -481 -501 -473 -497
rect -405 -501 -397 -497
rect -330 -501 -322 -497
rect -253 -501 -245 -497
rect -176 -501 -168 -497
rect -100 -501 -92 -497
rect -9 -501 -1 -497
rect 71 -500 79 -496
rect 150 -499 158 -495
rect 226 -498 234 -494
rect 540 -497 548 -493
rect 622 -497 630 -493
rect 1012 -492 1020 -488
rect 702 -497 710 -493
rect 831 -498 839 -494
rect 928 -498 936 -494
rect 1012 -500 1020 -496
rect -481 -526 -473 -522
rect -405 -526 -397 -522
rect -330 -526 -322 -522
rect -253 -526 -245 -522
rect -176 -526 -168 -522
rect -100 -526 -92 -522
rect -9 -526 -1 -522
rect 71 -525 79 -521
rect 150 -524 158 -520
rect 226 -523 234 -519
rect 540 -522 548 -518
rect 622 -522 630 -518
rect 702 -522 710 -518
rect 831 -523 839 -519
rect 928 -523 936 -519
rect -481 -534 -473 -530
rect -405 -534 -397 -530
rect -330 -534 -322 -530
rect -253 -534 -245 -530
rect -176 -534 -168 -530
rect -100 -534 -92 -530
rect -9 -534 -1 -530
rect 71 -533 79 -529
rect 150 -532 158 -528
rect 226 -531 234 -527
rect 540 -530 548 -526
rect 622 -530 630 -526
rect 1012 -525 1020 -521
rect 702 -530 710 -526
rect 831 -531 839 -527
rect 928 -531 936 -527
rect 1012 -533 1020 -529
rect -481 -549 -473 -545
rect -405 -549 -397 -545
rect -330 -549 -322 -545
rect -253 -549 -245 -545
rect -176 -549 -168 -545
rect -100 -549 -92 -545
rect -9 -549 -1 -545
rect 71 -548 79 -544
rect 150 -547 158 -543
rect 226 -546 234 -542
rect 540 -545 548 -541
rect 622 -545 630 -541
rect 702 -545 710 -541
rect 831 -546 839 -542
rect 928 -546 936 -542
rect -481 -557 -473 -553
rect -405 -557 -397 -553
rect -330 -557 -322 -553
rect -253 -557 -245 -553
rect -176 -557 -168 -553
rect -100 -557 -92 -553
rect -9 -557 -1 -553
rect 71 -556 79 -552
rect 150 -555 158 -551
rect 226 -554 234 -550
rect 540 -553 548 -549
rect 622 -553 630 -549
rect 1012 -548 1020 -544
rect 702 -553 710 -549
rect 831 -554 839 -550
rect 928 -554 936 -550
rect 1012 -556 1020 -552
rect 865 -632 869 -624
rect 873 -632 877 -624
rect 888 -632 892 -624
rect 896 -632 900 -624
rect 462 -658 466 -650
rect 470 -658 474 -650
rect 485 -658 489 -650
rect 493 -658 497 -650
rect 60 -678 64 -670
rect 68 -678 72 -670
rect 83 -678 87 -670
rect 91 -678 95 -670
rect 939 -662 943 -654
rect 947 -662 951 -654
rect 962 -662 966 -654
rect 970 -662 974 -654
rect 536 -688 540 -680
rect 544 -688 548 -680
rect 559 -688 563 -680
rect 567 -688 571 -680
rect 673 -686 677 -678
rect 681 -686 685 -678
rect 696 -686 700 -678
rect 704 -686 708 -678
rect 730 -686 734 -678
rect 738 -686 742 -678
rect 753 -686 757 -678
rect 761 -686 765 -678
rect 810 -684 814 -676
rect 818 -684 822 -676
rect 833 -684 837 -676
rect 841 -684 845 -676
rect 134 -708 138 -700
rect 142 -708 146 -700
rect 157 -708 161 -700
rect 165 -708 169 -700
rect -371 -716 -363 -712
rect -371 -724 -363 -720
rect -132 -732 -128 -724
rect -124 -732 -120 -724
rect -109 -732 -105 -724
rect -101 -732 -97 -724
rect -75 -732 -71 -724
rect -67 -732 -63 -724
rect -52 -732 -48 -724
rect -44 -732 -40 -724
rect 5 -730 9 -722
rect 13 -730 17 -722
rect 28 -730 32 -722
rect 36 -730 40 -722
rect -371 -739 -363 -735
rect -460 -744 -452 -740
rect -371 -747 -363 -743
rect -460 -752 -452 -748
rect 270 -712 274 -704
rect 278 -712 282 -704
rect 293 -712 297 -704
rect 301 -712 305 -704
rect 327 -712 331 -704
rect 335 -712 339 -704
rect 350 -712 354 -704
rect 358 -712 362 -704
rect 407 -710 411 -702
rect 415 -710 419 -702
rect 430 -710 434 -702
rect 438 -710 442 -702
rect 873 -707 877 -699
rect 881 -707 885 -699
rect 896 -707 900 -699
rect 904 -707 908 -699
rect 470 -733 474 -725
rect 478 -733 482 -725
rect 493 -733 497 -725
rect 501 -733 505 -725
rect 68 -753 72 -745
rect 76 -753 80 -745
rect 91 -753 95 -745
rect 99 -753 103 -745
rect -460 -767 -452 -763
rect -460 -775 -452 -771
rect -319 -771 -311 -767
rect -394 -779 -386 -775
rect -319 -779 -311 -775
rect -394 -787 -386 -783
rect -319 -794 -311 -790
rect -460 -801 -452 -797
rect -394 -802 -386 -798
rect -319 -802 -311 -798
rect -460 -809 -452 -805
rect -394 -810 -386 -806
rect -460 -824 -452 -820
rect -460 -832 -452 -828
rect -349 -845 -341 -841
rect -349 -853 -341 -849
rect -349 -868 -341 -864
rect -349 -876 -341 -872
rect -521 -927 -513 -923
rect -455 -927 -447 -923
rect -366 -928 -358 -924
rect -63 -927 -55 -923
rect -521 -935 -513 -931
rect -455 -935 -447 -931
rect -366 -936 -358 -932
rect -63 -935 -55 -931
rect -521 -950 -513 -946
rect -455 -950 -447 -946
rect -366 -951 -358 -947
rect -63 -950 -55 -946
rect 270 -946 278 -942
rect -521 -958 -513 -954
rect -455 -958 -447 -954
rect -366 -959 -358 -955
rect -152 -955 -144 -951
rect 270 -954 278 -950
rect -63 -958 -55 -954
rect -152 -963 -144 -959
rect 270 -969 278 -965
rect -152 -978 -144 -974
rect 181 -974 189 -970
rect 270 -977 278 -973
rect -455 -984 -447 -980
rect -314 -983 -306 -979
rect -152 -986 -144 -982
rect -11 -982 -3 -978
rect 181 -982 189 -978
rect -455 -992 -447 -988
rect -389 -991 -381 -987
rect -314 -991 -306 -987
rect -86 -990 -78 -986
rect 813 -985 821 -981
rect -11 -990 -3 -986
rect 813 -993 821 -989
rect -389 -999 -381 -995
rect -86 -998 -78 -994
rect 181 -997 189 -993
rect -534 -1008 -526 -1004
rect -455 -1007 -447 -1003
rect -314 -1006 -306 -1002
rect -11 -1005 -3 -1001
rect 181 -1005 189 -1001
rect 322 -1001 330 -997
rect -534 -1016 -526 -1012
rect -455 -1015 -447 -1011
rect -389 -1014 -381 -1010
rect -314 -1014 -306 -1010
rect -152 -1012 -144 -1008
rect -86 -1013 -78 -1009
rect -11 -1013 -3 -1009
rect 247 -1009 255 -1005
rect 322 -1009 330 -1005
rect 813 -1008 821 -1004
rect -389 -1022 -381 -1018
rect -152 -1020 -144 -1016
rect 247 -1017 255 -1013
rect 724 -1013 732 -1009
rect 813 -1016 821 -1012
rect -86 -1021 -78 -1017
rect 322 -1024 330 -1020
rect 724 -1021 732 -1017
rect -534 -1031 -526 -1027
rect -534 -1039 -526 -1035
rect -152 -1035 -144 -1031
rect 181 -1031 189 -1027
rect 247 -1032 255 -1028
rect 322 -1032 330 -1028
rect 181 -1039 189 -1035
rect -152 -1043 -144 -1039
rect 247 -1040 255 -1036
rect 724 -1036 732 -1032
rect 724 -1044 732 -1040
rect 865 -1040 873 -1036
rect -442 -1052 -434 -1048
rect 790 -1048 798 -1044
rect 865 -1048 873 -1044
rect -442 -1060 -434 -1056
rect -344 -1057 -336 -1053
rect -41 -1056 -33 -1052
rect 181 -1054 189 -1050
rect 790 -1056 798 -1052
rect -344 -1065 -336 -1061
rect -41 -1064 -33 -1060
rect 181 -1062 189 -1058
rect 865 -1063 873 -1059
rect 724 -1070 732 -1066
rect -442 -1075 -434 -1071
rect -442 -1083 -434 -1079
rect -344 -1080 -336 -1076
rect -41 -1079 -33 -1075
rect 292 -1075 300 -1071
rect 790 -1071 798 -1067
rect 865 -1071 873 -1067
rect 724 -1078 732 -1074
rect -344 -1088 -336 -1084
rect 790 -1079 798 -1075
rect 292 -1083 300 -1079
rect -41 -1087 -33 -1083
rect 724 -1093 732 -1089
rect 292 -1098 300 -1094
rect 724 -1101 732 -1097
rect 292 -1106 300 -1102
rect 835 -1114 843 -1110
rect 835 -1122 843 -1118
rect -213 -1138 -205 -1134
rect -147 -1138 -139 -1134
rect -58 -1139 -50 -1135
rect 835 -1137 843 -1133
rect -213 -1146 -205 -1142
rect -147 -1146 -139 -1142
rect -58 -1147 -50 -1143
rect 835 -1145 843 -1141
rect -213 -1161 -205 -1157
rect -147 -1161 -139 -1157
rect 120 -1157 128 -1153
rect 186 -1157 194 -1153
rect -58 -1162 -50 -1158
rect 275 -1158 283 -1154
rect -213 -1169 -205 -1165
rect 120 -1165 128 -1161
rect 186 -1165 194 -1161
rect -147 -1169 -139 -1165
rect 275 -1166 283 -1162
rect -58 -1170 -50 -1166
rect 120 -1180 128 -1176
rect 186 -1180 194 -1176
rect 275 -1181 283 -1177
rect 120 -1188 128 -1184
rect 186 -1188 194 -1184
rect 275 -1189 283 -1185
rect -147 -1195 -139 -1191
rect -6 -1194 2 -1190
rect 663 -1196 671 -1192
rect 729 -1196 737 -1192
rect -147 -1203 -139 -1199
rect -81 -1202 -73 -1198
rect -6 -1202 2 -1198
rect 818 -1197 826 -1193
rect 663 -1204 671 -1200
rect 729 -1204 737 -1200
rect 818 -1205 826 -1201
rect -81 -1210 -73 -1206
rect -226 -1219 -218 -1215
rect -147 -1218 -139 -1214
rect -6 -1217 2 -1213
rect 186 -1214 194 -1210
rect 327 -1213 335 -1209
rect -226 -1227 -218 -1223
rect -147 -1226 -139 -1222
rect -81 -1225 -73 -1221
rect -6 -1225 2 -1221
rect 186 -1222 194 -1218
rect 252 -1221 260 -1217
rect 327 -1221 335 -1217
rect 663 -1219 671 -1215
rect 729 -1219 737 -1215
rect 818 -1220 826 -1216
rect 252 -1229 260 -1225
rect 663 -1227 671 -1223
rect 729 -1227 737 -1223
rect 818 -1228 826 -1224
rect -81 -1233 -73 -1229
rect -226 -1242 -218 -1238
rect 107 -1238 115 -1234
rect 186 -1237 194 -1233
rect 327 -1236 335 -1232
rect 107 -1246 115 -1242
rect 186 -1245 194 -1241
rect 252 -1244 260 -1240
rect 327 -1244 335 -1240
rect -226 -1250 -218 -1246
rect 252 -1252 260 -1248
rect 729 -1253 737 -1249
rect 870 -1252 878 -1248
rect -134 -1263 -126 -1259
rect 107 -1261 115 -1257
rect 729 -1261 737 -1257
rect 795 -1260 803 -1256
rect 870 -1260 878 -1256
rect -134 -1271 -126 -1267
rect -36 -1268 -28 -1264
rect 107 -1269 115 -1265
rect 795 -1268 803 -1264
rect -36 -1276 -28 -1272
rect 650 -1277 658 -1273
rect 729 -1276 737 -1272
rect 870 -1275 878 -1271
rect -134 -1286 -126 -1282
rect 199 -1282 207 -1278
rect -134 -1294 -126 -1290
rect -36 -1291 -28 -1287
rect 199 -1290 207 -1286
rect 297 -1287 305 -1283
rect 650 -1285 658 -1281
rect 729 -1284 737 -1280
rect 795 -1283 803 -1279
rect 870 -1283 878 -1279
rect 795 -1291 803 -1287
rect 297 -1295 305 -1291
rect -36 -1299 -28 -1295
rect 650 -1300 658 -1296
rect 199 -1305 207 -1301
rect 199 -1313 207 -1309
rect 297 -1310 305 -1306
rect 650 -1308 658 -1304
rect 297 -1318 305 -1314
rect 742 -1321 750 -1317
rect 742 -1329 750 -1325
rect 840 -1326 848 -1322
rect 840 -1334 848 -1330
rect 742 -1344 750 -1340
rect 742 -1352 750 -1348
rect 840 -1349 848 -1345
rect 840 -1357 848 -1353
rect 516 -1508 524 -1504
rect 516 -1516 524 -1512
rect 516 -1531 524 -1527
rect 427 -1536 435 -1532
rect 516 -1539 524 -1535
rect 427 -1544 435 -1540
rect -127 -1556 -119 -1552
rect 427 -1559 435 -1555
rect -127 -1564 -119 -1560
rect 213 -1566 221 -1562
rect 427 -1567 435 -1563
rect 568 -1563 576 -1559
rect 213 -1574 221 -1570
rect 493 -1571 501 -1567
rect 568 -1571 576 -1567
rect -127 -1579 -119 -1575
rect 493 -1579 501 -1575
rect -216 -1584 -208 -1580
rect -127 -1587 -119 -1583
rect -216 -1592 -208 -1588
rect 213 -1589 221 -1585
rect 568 -1586 576 -1582
rect 124 -1594 132 -1590
rect 213 -1597 221 -1593
rect 427 -1593 435 -1589
rect 493 -1594 501 -1590
rect 568 -1594 576 -1590
rect 124 -1602 132 -1598
rect 427 -1601 435 -1597
rect 493 -1602 501 -1598
rect -216 -1607 -208 -1603
rect -432 -1612 -424 -1608
rect -216 -1615 -208 -1611
rect -75 -1611 -67 -1607
rect -432 -1620 -424 -1616
rect -150 -1619 -142 -1615
rect -75 -1619 -67 -1615
rect 124 -1617 132 -1613
rect 427 -1616 435 -1612
rect -150 -1627 -142 -1623
rect 124 -1625 132 -1621
rect 265 -1621 273 -1617
rect 427 -1624 435 -1620
rect 190 -1629 198 -1625
rect 265 -1629 273 -1625
rect -432 -1635 -424 -1631
rect -75 -1634 -67 -1630
rect -521 -1640 -513 -1636
rect 190 -1637 198 -1633
rect -432 -1643 -424 -1639
rect -216 -1641 -208 -1637
rect -150 -1642 -142 -1638
rect 538 -1637 546 -1633
rect -75 -1642 -67 -1638
rect -521 -1648 -513 -1644
rect 265 -1644 273 -1640
rect 538 -1645 546 -1641
rect -216 -1649 -208 -1645
rect -150 -1650 -142 -1646
rect 124 -1651 132 -1647
rect 190 -1652 198 -1648
rect 265 -1652 273 -1648
rect 124 -1659 132 -1655
rect -521 -1663 -513 -1659
rect 190 -1660 198 -1656
rect -521 -1671 -513 -1667
rect -380 -1667 -372 -1663
rect -216 -1664 -208 -1660
rect 538 -1660 546 -1656
rect -455 -1675 -447 -1671
rect -380 -1675 -372 -1671
rect 538 -1668 546 -1664
rect -216 -1672 -208 -1668
rect 124 -1674 132 -1670
rect -455 -1683 -447 -1679
rect -105 -1685 -97 -1681
rect 124 -1682 132 -1678
rect -380 -1690 -372 -1686
rect -105 -1693 -97 -1689
rect -521 -1697 -513 -1693
rect -455 -1698 -447 -1694
rect -380 -1698 -372 -1694
rect 235 -1695 243 -1691
rect -521 -1705 -513 -1701
rect -455 -1706 -447 -1702
rect 235 -1703 243 -1699
rect -105 -1708 -97 -1704
rect -105 -1716 -97 -1712
rect -521 -1720 -513 -1716
rect 235 -1718 243 -1714
rect 366 -1719 374 -1715
rect 432 -1719 440 -1715
rect -521 -1728 -513 -1724
rect 521 -1720 529 -1716
rect 235 -1726 243 -1722
rect 366 -1727 374 -1723
rect 432 -1727 440 -1723
rect 521 -1728 529 -1724
rect -410 -1741 -402 -1737
rect 366 -1742 374 -1738
rect 432 -1742 440 -1738
rect 521 -1743 529 -1739
rect -410 -1749 -402 -1745
rect 366 -1750 374 -1746
rect 432 -1750 440 -1746
rect 521 -1751 529 -1747
rect -410 -1764 -402 -1760
rect -277 -1767 -269 -1763
rect -211 -1767 -203 -1763
rect -410 -1772 -402 -1768
rect -122 -1768 -114 -1764
rect -277 -1775 -269 -1771
rect -211 -1775 -203 -1771
rect -122 -1776 -114 -1772
rect 63 -1777 71 -1773
rect 129 -1777 137 -1773
rect 218 -1778 226 -1774
rect 432 -1776 440 -1772
rect 573 -1775 581 -1771
rect 63 -1785 71 -1781
rect 129 -1785 137 -1781
rect 218 -1786 226 -1782
rect 432 -1784 440 -1780
rect 498 -1783 506 -1779
rect 573 -1783 581 -1779
rect -277 -1790 -269 -1786
rect -211 -1790 -203 -1786
rect -122 -1791 -114 -1787
rect 498 -1791 506 -1787
rect -277 -1798 -269 -1794
rect -211 -1798 -203 -1794
rect -122 -1799 -114 -1795
rect 63 -1800 71 -1796
rect 129 -1800 137 -1796
rect 218 -1801 226 -1797
rect 353 -1800 361 -1796
rect 432 -1799 440 -1795
rect 573 -1798 581 -1794
rect 63 -1808 71 -1804
rect 129 -1808 137 -1804
rect 218 -1809 226 -1805
rect 353 -1808 361 -1804
rect 432 -1807 440 -1803
rect 498 -1806 506 -1802
rect 573 -1806 581 -1802
rect 498 -1814 506 -1810
rect -582 -1823 -574 -1819
rect -516 -1823 -508 -1819
rect -427 -1824 -419 -1820
rect -211 -1824 -203 -1820
rect -70 -1823 -62 -1819
rect 353 -1823 361 -1819
rect -582 -1831 -574 -1827
rect -516 -1831 -508 -1827
rect -427 -1832 -419 -1828
rect -211 -1832 -203 -1828
rect -145 -1831 -137 -1827
rect -70 -1831 -62 -1827
rect 129 -1834 137 -1830
rect 270 -1833 278 -1829
rect 353 -1831 361 -1827
rect -145 -1839 -137 -1835
rect 129 -1842 137 -1838
rect 195 -1841 203 -1837
rect 270 -1841 278 -1837
rect -582 -1846 -574 -1842
rect -516 -1846 -508 -1842
rect -427 -1847 -419 -1843
rect -582 -1854 -574 -1850
rect -290 -1848 -282 -1844
rect -211 -1847 -203 -1843
rect -70 -1846 -62 -1842
rect -516 -1854 -508 -1850
rect 445 -1844 453 -1840
rect 195 -1849 203 -1845
rect -427 -1855 -419 -1851
rect -290 -1856 -282 -1852
rect -211 -1855 -203 -1851
rect -145 -1854 -137 -1850
rect -70 -1854 -62 -1850
rect 445 -1852 453 -1848
rect 543 -1849 551 -1845
rect -145 -1862 -137 -1858
rect 50 -1858 58 -1854
rect 129 -1857 137 -1853
rect 270 -1856 278 -1852
rect 543 -1857 551 -1853
rect 50 -1866 58 -1862
rect 129 -1865 137 -1861
rect 195 -1864 203 -1860
rect 270 -1864 278 -1860
rect -290 -1871 -282 -1867
rect 445 -1867 453 -1863
rect 195 -1872 203 -1868
rect -516 -1880 -508 -1876
rect -375 -1879 -367 -1875
rect 445 -1875 453 -1871
rect 543 -1872 551 -1868
rect -290 -1879 -282 -1875
rect 50 -1881 58 -1877
rect 543 -1880 551 -1876
rect -516 -1888 -508 -1884
rect -450 -1887 -442 -1883
rect -375 -1887 -367 -1883
rect -450 -1895 -442 -1891
rect -198 -1892 -190 -1888
rect 50 -1889 58 -1885
rect -595 -1904 -587 -1900
rect -516 -1903 -508 -1899
rect -375 -1902 -367 -1898
rect -198 -1900 -190 -1896
rect -100 -1897 -92 -1893
rect -100 -1905 -92 -1901
rect 142 -1902 150 -1898
rect -595 -1912 -587 -1908
rect -516 -1911 -508 -1907
rect -450 -1910 -442 -1906
rect -375 -1910 -367 -1906
rect 142 -1910 150 -1906
rect 240 -1907 248 -1903
rect -450 -1918 -442 -1914
rect -198 -1915 -190 -1911
rect 240 -1915 248 -1911
rect -198 -1923 -190 -1919
rect -100 -1920 -92 -1916
rect -595 -1927 -587 -1923
rect -100 -1928 -92 -1924
rect 142 -1925 150 -1921
rect -595 -1935 -587 -1931
rect 142 -1933 150 -1929
rect 240 -1930 248 -1926
rect 240 -1938 248 -1934
rect -503 -1948 -495 -1944
rect -503 -1956 -495 -1952
rect -405 -1953 -397 -1949
rect -405 -1961 -397 -1957
rect -503 -1971 -495 -1967
rect -503 -1979 -495 -1975
rect -405 -1976 -397 -1972
rect -405 -1984 -397 -1980
rect 446 -2047 450 -2039
rect 454 -2047 458 -2039
rect 469 -2047 473 -2039
rect 477 -2047 481 -2039
rect 520 -2077 524 -2069
rect 528 -2077 532 -2069
rect 543 -2077 547 -2069
rect 551 -2077 555 -2069
rect 254 -2101 258 -2093
rect 262 -2101 266 -2093
rect 277 -2101 281 -2093
rect 285 -2101 289 -2093
rect 311 -2101 315 -2093
rect 319 -2101 323 -2093
rect 334 -2101 338 -2093
rect 342 -2101 346 -2093
rect 391 -2099 395 -2091
rect 399 -2099 403 -2091
rect 414 -2099 418 -2091
rect 422 -2099 426 -2091
rect 454 -2122 458 -2114
rect 462 -2122 466 -2114
rect 477 -2122 481 -2114
rect 485 -2122 489 -2114
<< polysilicon >>
rect -517 -473 -513 -471
rect -507 -473 -481 -471
rect -473 -473 -470 -471
rect -441 -473 -437 -471
rect -431 -473 -405 -471
rect -397 -473 -394 -471
rect -366 -473 -362 -471
rect -356 -473 -330 -471
rect -322 -473 -319 -471
rect -289 -473 -285 -471
rect -279 -473 -253 -471
rect -245 -473 -242 -471
rect -212 -473 -208 -471
rect -202 -473 -176 -471
rect -168 -473 -165 -471
rect -136 -473 -132 -471
rect -126 -473 -100 -471
rect -92 -473 -89 -471
rect -45 -473 -41 -471
rect -35 -473 -9 -471
rect -1 -473 2 -471
rect 35 -472 39 -470
rect 45 -472 71 -470
rect 79 -472 82 -470
rect 114 -471 118 -469
rect 124 -471 150 -469
rect 158 -471 161 -469
rect 190 -470 194 -468
rect 200 -470 226 -468
rect 234 -470 237 -468
rect 504 -469 508 -467
rect 514 -469 540 -467
rect 548 -469 551 -467
rect 586 -469 590 -467
rect 596 -469 622 -467
rect 630 -469 633 -467
rect 666 -469 670 -467
rect 676 -469 702 -467
rect 710 -469 713 -467
rect 795 -470 799 -468
rect 805 -470 831 -468
rect 839 -470 842 -468
rect 892 -470 896 -468
rect 902 -470 928 -468
rect 936 -470 939 -468
rect 976 -472 980 -470
rect 986 -472 1012 -470
rect 1020 -472 1023 -470
rect -517 -496 -513 -494
rect -507 -496 -481 -494
rect -473 -496 -470 -494
rect -441 -496 -437 -494
rect -431 -496 -405 -494
rect -397 -496 -394 -494
rect -366 -496 -362 -494
rect -356 -496 -330 -494
rect -322 -496 -319 -494
rect -289 -496 -285 -494
rect -279 -496 -253 -494
rect -245 -496 -242 -494
rect -212 -496 -208 -494
rect -202 -496 -176 -494
rect -168 -496 -165 -494
rect -136 -496 -132 -494
rect -126 -496 -100 -494
rect -92 -496 -89 -494
rect -45 -496 -41 -494
rect -35 -496 -9 -494
rect -1 -496 2 -494
rect 35 -495 39 -493
rect 45 -495 71 -493
rect 79 -495 82 -493
rect 114 -494 118 -492
rect 124 -494 150 -492
rect 158 -494 161 -492
rect 190 -493 194 -491
rect 200 -493 226 -491
rect 234 -493 237 -491
rect 504 -492 508 -490
rect 514 -492 540 -490
rect 548 -492 551 -490
rect 586 -492 590 -490
rect 596 -492 622 -490
rect 630 -492 633 -490
rect 666 -492 670 -490
rect 676 -492 702 -490
rect 710 -492 713 -490
rect 795 -493 799 -491
rect 805 -493 831 -491
rect 839 -493 842 -491
rect 892 -493 896 -491
rect 902 -493 928 -491
rect 936 -493 939 -491
rect 976 -495 980 -493
rect 986 -495 1012 -493
rect 1020 -495 1023 -493
rect -517 -529 -513 -527
rect -507 -529 -481 -527
rect -473 -529 -470 -527
rect -441 -529 -437 -527
rect -431 -529 -405 -527
rect -397 -529 -394 -527
rect -366 -529 -362 -527
rect -356 -529 -330 -527
rect -322 -529 -319 -527
rect -289 -529 -285 -527
rect -279 -529 -253 -527
rect -245 -529 -242 -527
rect -212 -529 -208 -527
rect -202 -529 -176 -527
rect -168 -529 -165 -527
rect -136 -529 -132 -527
rect -126 -529 -100 -527
rect -92 -529 -89 -527
rect -45 -529 -41 -527
rect -35 -529 -9 -527
rect -1 -529 2 -527
rect 35 -528 39 -526
rect 45 -528 71 -526
rect 79 -528 82 -526
rect 114 -527 118 -525
rect 124 -527 150 -525
rect 158 -527 161 -525
rect 190 -526 194 -524
rect 200 -526 226 -524
rect 234 -526 237 -524
rect 504 -525 508 -523
rect 514 -525 540 -523
rect 548 -525 551 -523
rect 586 -525 590 -523
rect 596 -525 622 -523
rect 630 -525 633 -523
rect 666 -525 670 -523
rect 676 -525 702 -523
rect 710 -525 713 -523
rect 795 -526 799 -524
rect 805 -526 831 -524
rect 839 -526 842 -524
rect 892 -526 896 -524
rect 902 -526 928 -524
rect 936 -526 939 -524
rect 976 -528 980 -526
rect 986 -528 1012 -526
rect 1020 -528 1023 -526
rect -517 -552 -513 -550
rect -507 -552 -481 -550
rect -473 -552 -470 -550
rect -441 -552 -437 -550
rect -431 -552 -405 -550
rect -397 -552 -394 -550
rect -366 -552 -362 -550
rect -356 -552 -330 -550
rect -322 -552 -319 -550
rect -289 -552 -285 -550
rect -279 -552 -253 -550
rect -245 -552 -242 -550
rect -212 -552 -208 -550
rect -202 -552 -176 -550
rect -168 -552 -165 -550
rect -136 -552 -132 -550
rect -126 -552 -100 -550
rect -92 -552 -89 -550
rect -45 -552 -41 -550
rect -35 -552 -9 -550
rect -1 -552 2 -550
rect 35 -551 39 -549
rect 45 -551 71 -549
rect 79 -551 82 -549
rect 114 -550 118 -548
rect 124 -550 150 -548
rect 158 -550 161 -548
rect 190 -549 194 -547
rect 200 -549 226 -547
rect 234 -549 237 -547
rect 504 -548 508 -546
rect 514 -548 540 -546
rect 548 -548 551 -546
rect 586 -548 590 -546
rect 596 -548 622 -546
rect 630 -548 633 -546
rect 666 -548 670 -546
rect 676 -548 702 -546
rect 710 -548 713 -546
rect 795 -549 799 -547
rect 805 -549 831 -547
rect 839 -549 842 -547
rect 892 -549 896 -547
rect 902 -549 928 -547
rect 936 -549 939 -547
rect 976 -551 980 -549
rect 986 -551 1012 -549
rect 1020 -551 1023 -549
rect 870 -624 872 -621
rect 893 -624 895 -621
rect 467 -650 469 -647
rect 490 -650 492 -647
rect 870 -658 872 -632
rect 893 -658 895 -632
rect 944 -654 946 -651
rect 967 -654 969 -651
rect 65 -670 67 -667
rect 88 -670 90 -667
rect 65 -704 67 -678
rect 88 -704 90 -678
rect 467 -684 469 -658
rect 490 -684 492 -658
rect 870 -668 872 -664
rect 893 -668 895 -664
rect 541 -680 543 -677
rect 564 -680 566 -677
rect 678 -678 680 -675
rect 701 -678 703 -675
rect 735 -678 737 -675
rect 758 -678 760 -675
rect 815 -676 817 -673
rect 838 -676 840 -673
rect 467 -694 469 -690
rect 490 -694 492 -690
rect 139 -700 141 -697
rect 162 -700 164 -697
rect 275 -704 277 -701
rect 298 -704 300 -701
rect 332 -704 334 -701
rect 355 -704 357 -701
rect 412 -702 414 -699
rect 435 -702 437 -699
rect 65 -714 67 -710
rect 88 -714 90 -710
rect -407 -719 -403 -717
rect -397 -719 -371 -717
rect -363 -719 -360 -717
rect -127 -724 -125 -721
rect -104 -724 -102 -721
rect -70 -724 -68 -721
rect -47 -724 -45 -721
rect 10 -722 12 -719
rect 33 -722 35 -719
rect -407 -742 -403 -740
rect -397 -742 -371 -740
rect -363 -742 -360 -740
rect -496 -747 -492 -745
rect -486 -747 -460 -745
rect -452 -747 -449 -745
rect -127 -758 -125 -732
rect -104 -758 -102 -732
rect -70 -758 -68 -732
rect -47 -758 -45 -732
rect 10 -756 12 -730
rect 33 -756 35 -730
rect 139 -734 141 -708
rect 162 -734 164 -708
rect 275 -738 277 -712
rect 298 -738 300 -712
rect 332 -738 334 -712
rect 355 -738 357 -712
rect 412 -736 414 -710
rect 435 -736 437 -710
rect 541 -714 543 -688
rect 564 -714 566 -688
rect 678 -712 680 -686
rect 701 -712 703 -686
rect 735 -712 737 -686
rect 758 -712 760 -686
rect 815 -710 817 -684
rect 838 -710 840 -684
rect 944 -688 946 -662
rect 967 -688 969 -662
rect 878 -699 880 -696
rect 901 -699 903 -696
rect 944 -698 946 -694
rect 967 -698 969 -694
rect 475 -725 477 -722
rect 498 -725 500 -722
rect 541 -724 543 -720
rect 564 -724 566 -720
rect 678 -722 680 -718
rect 701 -722 703 -718
rect 735 -722 737 -718
rect 758 -722 760 -718
rect 815 -720 817 -716
rect 838 -720 840 -716
rect 878 -733 880 -707
rect 901 -733 903 -707
rect 73 -745 75 -742
rect 96 -745 98 -742
rect 139 -744 141 -740
rect 162 -744 164 -740
rect 275 -748 277 -744
rect 298 -748 300 -744
rect 332 -748 334 -744
rect 355 -748 357 -744
rect 412 -746 414 -742
rect 435 -746 437 -742
rect -496 -770 -492 -768
rect -486 -770 -460 -768
rect -452 -770 -449 -768
rect -127 -768 -125 -764
rect -104 -768 -102 -764
rect -70 -768 -68 -764
rect -47 -768 -45 -764
rect 10 -766 12 -762
rect 33 -766 35 -762
rect -355 -774 -351 -772
rect -345 -774 -319 -772
rect -311 -774 -308 -772
rect 73 -779 75 -753
rect 96 -779 98 -753
rect 475 -759 477 -733
rect 498 -759 500 -733
rect 878 -743 880 -739
rect 901 -743 903 -739
rect 475 -769 477 -765
rect 498 -769 500 -765
rect -430 -782 -426 -780
rect -420 -782 -394 -780
rect -386 -782 -383 -780
rect 73 -789 75 -785
rect 96 -789 98 -785
rect -355 -797 -351 -795
rect -345 -797 -319 -795
rect -311 -797 -308 -795
rect -496 -804 -492 -802
rect -486 -804 -460 -802
rect -452 -804 -449 -802
rect -430 -805 -426 -803
rect -420 -805 -394 -803
rect -386 -805 -383 -803
rect -496 -827 -492 -825
rect -486 -827 -460 -825
rect -452 -827 -449 -825
rect -385 -848 -381 -846
rect -375 -848 -349 -846
rect -341 -848 -338 -846
rect -385 -871 -381 -869
rect -375 -871 -349 -869
rect -341 -871 -338 -869
rect -557 -930 -553 -928
rect -547 -930 -521 -928
rect -513 -930 -510 -928
rect -491 -930 -487 -928
rect -481 -930 -455 -928
rect -447 -930 -444 -928
rect -402 -931 -398 -929
rect -392 -931 -366 -929
rect -358 -931 -355 -929
rect -99 -930 -95 -928
rect -89 -930 -63 -928
rect -55 -930 -52 -928
rect -557 -953 -553 -951
rect -547 -953 -521 -951
rect -513 -953 -510 -951
rect -491 -953 -487 -951
rect -481 -953 -455 -951
rect -447 -953 -444 -951
rect 234 -949 238 -947
rect 244 -949 270 -947
rect 278 -949 281 -947
rect -402 -954 -398 -952
rect -392 -954 -366 -952
rect -358 -954 -355 -952
rect -99 -953 -95 -951
rect -89 -953 -63 -951
rect -55 -953 -52 -951
rect -188 -958 -184 -956
rect -178 -958 -152 -956
rect -144 -958 -141 -956
rect 234 -972 238 -970
rect 244 -972 270 -970
rect 278 -972 281 -970
rect 145 -977 149 -975
rect 155 -977 181 -975
rect 189 -977 192 -975
rect -188 -981 -184 -979
rect -178 -981 -152 -979
rect -144 -981 -141 -979
rect -491 -987 -487 -985
rect -481 -987 -455 -985
rect -447 -987 -444 -985
rect -350 -986 -346 -984
rect -340 -986 -314 -984
rect -306 -986 -303 -984
rect -47 -985 -43 -983
rect -37 -985 -11 -983
rect -3 -985 0 -983
rect 777 -988 781 -986
rect 787 -988 813 -986
rect 821 -988 824 -986
rect -425 -994 -421 -992
rect -415 -994 -389 -992
rect -381 -994 -378 -992
rect -122 -993 -118 -991
rect -112 -993 -86 -991
rect -78 -993 -75 -991
rect 145 -1000 149 -998
rect 155 -1000 181 -998
rect 189 -1000 192 -998
rect 286 -1004 290 -1002
rect 296 -1004 322 -1002
rect 330 -1004 333 -1002
rect -570 -1011 -566 -1009
rect -560 -1011 -534 -1009
rect -526 -1011 -523 -1009
rect -491 -1010 -487 -1008
rect -481 -1010 -455 -1008
rect -447 -1010 -444 -1008
rect -350 -1009 -346 -1007
rect -340 -1009 -314 -1007
rect -306 -1009 -303 -1007
rect -47 -1008 -43 -1006
rect -37 -1008 -11 -1006
rect -3 -1008 0 -1006
rect -188 -1015 -184 -1013
rect -178 -1015 -152 -1013
rect -144 -1015 -141 -1013
rect 211 -1012 215 -1010
rect 221 -1012 247 -1010
rect 255 -1012 258 -1010
rect -425 -1017 -421 -1015
rect -415 -1017 -389 -1015
rect -381 -1017 -378 -1015
rect -122 -1016 -118 -1014
rect -112 -1016 -86 -1014
rect -78 -1016 -75 -1014
rect 777 -1011 781 -1009
rect 787 -1011 813 -1009
rect 821 -1011 824 -1009
rect 688 -1016 692 -1014
rect 698 -1016 724 -1014
rect 732 -1016 735 -1014
rect 286 -1027 290 -1025
rect 296 -1027 322 -1025
rect 330 -1027 333 -1025
rect -570 -1034 -566 -1032
rect -560 -1034 -534 -1032
rect -526 -1034 -523 -1032
rect 145 -1034 149 -1032
rect 155 -1034 181 -1032
rect 189 -1034 192 -1032
rect -188 -1038 -184 -1036
rect -178 -1038 -152 -1036
rect -144 -1038 -141 -1036
rect 211 -1035 215 -1033
rect 221 -1035 247 -1033
rect 255 -1035 258 -1033
rect 688 -1039 692 -1037
rect 698 -1039 724 -1037
rect 732 -1039 735 -1037
rect 829 -1043 833 -1041
rect 839 -1043 865 -1041
rect 873 -1043 876 -1041
rect -478 -1055 -474 -1053
rect -468 -1055 -442 -1053
rect -434 -1055 -431 -1053
rect 754 -1051 758 -1049
rect 764 -1051 790 -1049
rect 798 -1051 801 -1049
rect 145 -1057 149 -1055
rect 155 -1057 181 -1055
rect 189 -1057 192 -1055
rect -380 -1060 -376 -1058
rect -370 -1060 -344 -1058
rect -336 -1060 -333 -1058
rect -77 -1059 -73 -1057
rect -67 -1059 -41 -1057
rect -33 -1059 -30 -1057
rect 829 -1066 833 -1064
rect 839 -1066 865 -1064
rect 873 -1066 876 -1064
rect -478 -1078 -474 -1076
rect -468 -1078 -442 -1076
rect -434 -1078 -431 -1076
rect 688 -1073 692 -1071
rect 698 -1073 724 -1071
rect 732 -1073 735 -1071
rect 256 -1078 260 -1076
rect 266 -1078 292 -1076
rect 300 -1078 303 -1076
rect 754 -1074 758 -1072
rect 764 -1074 790 -1072
rect 798 -1074 801 -1072
rect -380 -1083 -376 -1081
rect -370 -1083 -344 -1081
rect -336 -1083 -333 -1081
rect -77 -1082 -73 -1080
rect -67 -1082 -41 -1080
rect -33 -1082 -30 -1080
rect 688 -1096 692 -1094
rect 698 -1096 724 -1094
rect 732 -1096 735 -1094
rect 256 -1101 260 -1099
rect 266 -1101 292 -1099
rect 300 -1101 303 -1099
rect 799 -1117 803 -1115
rect 809 -1117 835 -1115
rect 843 -1117 846 -1115
rect -249 -1141 -245 -1139
rect -239 -1141 -213 -1139
rect -205 -1141 -202 -1139
rect -183 -1141 -179 -1139
rect -173 -1141 -147 -1139
rect -139 -1141 -136 -1139
rect 799 -1140 803 -1138
rect 809 -1140 835 -1138
rect 843 -1140 846 -1138
rect -94 -1142 -90 -1140
rect -84 -1142 -58 -1140
rect -50 -1142 -47 -1140
rect -249 -1164 -245 -1162
rect -239 -1164 -213 -1162
rect -205 -1164 -202 -1162
rect -183 -1164 -179 -1162
rect -173 -1164 -147 -1162
rect -139 -1164 -136 -1162
rect 84 -1160 88 -1158
rect 94 -1160 120 -1158
rect 128 -1160 131 -1158
rect 150 -1160 154 -1158
rect 160 -1160 186 -1158
rect 194 -1160 197 -1158
rect -94 -1165 -90 -1163
rect -84 -1165 -58 -1163
rect -50 -1165 -47 -1163
rect 239 -1161 243 -1159
rect 249 -1161 275 -1159
rect 283 -1161 286 -1159
rect 84 -1183 88 -1181
rect 94 -1183 120 -1181
rect 128 -1183 131 -1181
rect 150 -1183 154 -1181
rect 160 -1183 186 -1181
rect 194 -1183 197 -1181
rect 239 -1184 243 -1182
rect 249 -1184 275 -1182
rect 283 -1184 286 -1182
rect -183 -1198 -179 -1196
rect -173 -1198 -147 -1196
rect -139 -1198 -136 -1196
rect -42 -1197 -38 -1195
rect -32 -1197 -6 -1195
rect 2 -1197 5 -1195
rect 627 -1199 631 -1197
rect 637 -1199 663 -1197
rect 671 -1199 674 -1197
rect 693 -1199 697 -1197
rect 703 -1199 729 -1197
rect 737 -1199 740 -1197
rect -117 -1205 -113 -1203
rect -107 -1205 -81 -1203
rect -73 -1205 -70 -1203
rect 782 -1200 786 -1198
rect 792 -1200 818 -1198
rect 826 -1200 829 -1198
rect 150 -1217 154 -1215
rect 160 -1217 186 -1215
rect 194 -1217 197 -1215
rect 291 -1216 295 -1214
rect 301 -1216 327 -1214
rect 335 -1216 338 -1214
rect -262 -1222 -258 -1220
rect -252 -1222 -226 -1220
rect -218 -1222 -215 -1220
rect -183 -1221 -179 -1219
rect -173 -1221 -147 -1219
rect -139 -1221 -136 -1219
rect -42 -1220 -38 -1218
rect -32 -1220 -6 -1218
rect 2 -1220 5 -1218
rect 627 -1222 631 -1220
rect 637 -1222 663 -1220
rect 671 -1222 674 -1220
rect 693 -1222 697 -1220
rect 703 -1222 729 -1220
rect 737 -1222 740 -1220
rect 216 -1224 220 -1222
rect 226 -1224 252 -1222
rect 260 -1224 263 -1222
rect -117 -1228 -113 -1226
rect -107 -1228 -81 -1226
rect -73 -1228 -70 -1226
rect 782 -1223 786 -1221
rect 792 -1223 818 -1221
rect 826 -1223 829 -1221
rect 71 -1241 75 -1239
rect 81 -1241 107 -1239
rect 115 -1241 118 -1239
rect 150 -1240 154 -1238
rect 160 -1240 186 -1238
rect 194 -1240 197 -1238
rect 291 -1239 295 -1237
rect 301 -1239 327 -1237
rect 335 -1239 338 -1237
rect -262 -1245 -258 -1243
rect -252 -1245 -226 -1243
rect -218 -1245 -215 -1243
rect 216 -1247 220 -1245
rect 226 -1247 252 -1245
rect 260 -1247 263 -1245
rect 693 -1256 697 -1254
rect 703 -1256 729 -1254
rect 737 -1256 740 -1254
rect 834 -1255 838 -1253
rect 844 -1255 870 -1253
rect 878 -1255 881 -1253
rect 71 -1264 75 -1262
rect 81 -1264 107 -1262
rect 115 -1264 118 -1262
rect 759 -1263 763 -1261
rect 769 -1263 795 -1261
rect 803 -1263 806 -1261
rect -170 -1266 -166 -1264
rect -160 -1266 -134 -1264
rect -126 -1266 -123 -1264
rect -72 -1271 -68 -1269
rect -62 -1271 -36 -1269
rect -28 -1271 -25 -1269
rect 614 -1280 618 -1278
rect 624 -1280 650 -1278
rect 658 -1280 661 -1278
rect 693 -1279 697 -1277
rect 703 -1279 729 -1277
rect 737 -1279 740 -1277
rect 834 -1278 838 -1276
rect 844 -1278 870 -1276
rect 878 -1278 881 -1276
rect 163 -1285 167 -1283
rect 173 -1285 199 -1283
rect 207 -1285 210 -1283
rect -170 -1289 -166 -1287
rect -160 -1289 -134 -1287
rect -126 -1289 -123 -1287
rect 759 -1286 763 -1284
rect 769 -1286 795 -1284
rect 803 -1286 806 -1284
rect 261 -1290 265 -1288
rect 271 -1290 297 -1288
rect 305 -1290 308 -1288
rect -72 -1294 -68 -1292
rect -62 -1294 -36 -1292
rect -28 -1294 -25 -1292
rect 614 -1303 618 -1301
rect 624 -1303 650 -1301
rect 658 -1303 661 -1301
rect 163 -1308 167 -1306
rect 173 -1308 199 -1306
rect 207 -1308 210 -1306
rect 261 -1313 265 -1311
rect 271 -1313 297 -1311
rect 305 -1313 308 -1311
rect 706 -1324 710 -1322
rect 716 -1324 742 -1322
rect 750 -1324 753 -1322
rect 804 -1329 808 -1327
rect 814 -1329 840 -1327
rect 848 -1329 851 -1327
rect 706 -1347 710 -1345
rect 716 -1347 742 -1345
rect 750 -1347 753 -1345
rect 804 -1352 808 -1350
rect 814 -1352 840 -1350
rect 848 -1352 851 -1350
rect 480 -1511 484 -1509
rect 490 -1511 516 -1509
rect 524 -1511 527 -1509
rect 480 -1534 484 -1532
rect 490 -1534 516 -1532
rect 524 -1534 527 -1532
rect 391 -1539 395 -1537
rect 401 -1539 427 -1537
rect 435 -1539 438 -1537
rect -163 -1559 -159 -1557
rect -153 -1559 -127 -1557
rect -119 -1559 -116 -1557
rect 391 -1562 395 -1560
rect 401 -1562 427 -1560
rect 435 -1562 438 -1560
rect 532 -1566 536 -1564
rect 542 -1566 568 -1564
rect 576 -1566 579 -1564
rect 177 -1569 181 -1567
rect 187 -1569 213 -1567
rect 221 -1569 224 -1567
rect 457 -1574 461 -1572
rect 467 -1574 493 -1572
rect 501 -1574 504 -1572
rect -163 -1582 -159 -1580
rect -153 -1582 -127 -1580
rect -119 -1582 -116 -1580
rect -252 -1587 -248 -1585
rect -242 -1587 -216 -1585
rect -208 -1587 -205 -1585
rect 532 -1589 536 -1587
rect 542 -1589 568 -1587
rect 576 -1589 579 -1587
rect 177 -1592 181 -1590
rect 187 -1592 213 -1590
rect 221 -1592 224 -1590
rect 88 -1597 92 -1595
rect 98 -1597 124 -1595
rect 132 -1597 135 -1595
rect 391 -1596 395 -1594
rect 401 -1596 427 -1594
rect 435 -1596 438 -1594
rect 457 -1597 461 -1595
rect 467 -1597 493 -1595
rect 501 -1597 504 -1595
rect -252 -1610 -248 -1608
rect -242 -1610 -216 -1608
rect -208 -1610 -205 -1608
rect -468 -1615 -464 -1613
rect -458 -1615 -432 -1613
rect -424 -1615 -421 -1613
rect -111 -1614 -107 -1612
rect -101 -1614 -75 -1612
rect -67 -1614 -64 -1612
rect 88 -1620 92 -1618
rect 98 -1620 124 -1618
rect 132 -1620 135 -1618
rect -186 -1622 -182 -1620
rect -176 -1622 -150 -1620
rect -142 -1622 -139 -1620
rect 391 -1619 395 -1617
rect 401 -1619 427 -1617
rect 435 -1619 438 -1617
rect 229 -1624 233 -1622
rect 239 -1624 265 -1622
rect 273 -1624 276 -1622
rect 154 -1632 158 -1630
rect 164 -1632 190 -1630
rect 198 -1632 201 -1630
rect -468 -1638 -464 -1636
rect -458 -1638 -432 -1636
rect -424 -1638 -421 -1636
rect -111 -1637 -107 -1635
rect -101 -1637 -75 -1635
rect -67 -1637 -64 -1635
rect -557 -1643 -553 -1641
rect -547 -1643 -521 -1641
rect -513 -1643 -510 -1641
rect -252 -1644 -248 -1642
rect -242 -1644 -216 -1642
rect -208 -1644 -205 -1642
rect 502 -1640 506 -1638
rect 512 -1640 538 -1638
rect 546 -1640 549 -1638
rect -186 -1645 -182 -1643
rect -176 -1645 -150 -1643
rect -142 -1645 -139 -1643
rect 229 -1647 233 -1645
rect 239 -1647 265 -1645
rect 273 -1647 276 -1645
rect 88 -1654 92 -1652
rect 98 -1654 124 -1652
rect 132 -1654 135 -1652
rect 154 -1655 158 -1653
rect 164 -1655 190 -1653
rect 198 -1655 201 -1653
rect -557 -1666 -553 -1664
rect -547 -1666 -521 -1664
rect -513 -1666 -510 -1664
rect 502 -1663 506 -1661
rect 512 -1663 538 -1661
rect 546 -1663 549 -1661
rect -252 -1667 -248 -1665
rect -242 -1667 -216 -1665
rect -208 -1667 -205 -1665
rect -416 -1670 -412 -1668
rect -406 -1670 -380 -1668
rect -372 -1670 -369 -1668
rect -491 -1678 -487 -1676
rect -481 -1678 -455 -1676
rect -447 -1678 -444 -1676
rect 88 -1677 92 -1675
rect 98 -1677 124 -1675
rect 132 -1677 135 -1675
rect -141 -1688 -137 -1686
rect -131 -1688 -105 -1686
rect -97 -1688 -94 -1686
rect -416 -1693 -412 -1691
rect -406 -1693 -380 -1691
rect -372 -1693 -369 -1691
rect -557 -1700 -553 -1698
rect -547 -1700 -521 -1698
rect -513 -1700 -510 -1698
rect 199 -1698 203 -1696
rect 209 -1698 235 -1696
rect 243 -1698 246 -1696
rect -491 -1701 -487 -1699
rect -481 -1701 -455 -1699
rect -447 -1701 -444 -1699
rect -141 -1711 -137 -1709
rect -131 -1711 -105 -1709
rect -97 -1711 -94 -1709
rect 199 -1721 203 -1719
rect 209 -1721 235 -1719
rect 243 -1721 246 -1719
rect -557 -1723 -553 -1721
rect -547 -1723 -521 -1721
rect -513 -1723 -510 -1721
rect 330 -1722 334 -1720
rect 340 -1722 366 -1720
rect 374 -1722 377 -1720
rect 396 -1722 400 -1720
rect 406 -1722 432 -1720
rect 440 -1722 443 -1720
rect 485 -1723 489 -1721
rect 495 -1723 521 -1721
rect 529 -1723 532 -1721
rect -446 -1744 -442 -1742
rect -436 -1744 -410 -1742
rect -402 -1744 -399 -1742
rect 330 -1745 334 -1743
rect 340 -1745 366 -1743
rect 374 -1745 377 -1743
rect 396 -1745 400 -1743
rect 406 -1745 432 -1743
rect 440 -1745 443 -1743
rect 485 -1746 489 -1744
rect 495 -1746 521 -1744
rect 529 -1746 532 -1744
rect -446 -1767 -442 -1765
rect -436 -1767 -410 -1765
rect -402 -1767 -399 -1765
rect -313 -1770 -309 -1768
rect -303 -1770 -277 -1768
rect -269 -1770 -266 -1768
rect -247 -1770 -243 -1768
rect -237 -1770 -211 -1768
rect -203 -1770 -200 -1768
rect -158 -1771 -154 -1769
rect -148 -1771 -122 -1769
rect -114 -1771 -111 -1769
rect 27 -1780 31 -1778
rect 37 -1780 63 -1778
rect 71 -1780 74 -1778
rect 93 -1780 97 -1778
rect 103 -1780 129 -1778
rect 137 -1780 140 -1778
rect 396 -1779 400 -1777
rect 406 -1779 432 -1777
rect 440 -1779 443 -1777
rect 537 -1778 541 -1776
rect 547 -1778 573 -1776
rect 581 -1778 584 -1776
rect 182 -1781 186 -1779
rect 192 -1781 218 -1779
rect 226 -1781 229 -1779
rect 462 -1786 466 -1784
rect 472 -1786 498 -1784
rect 506 -1786 509 -1784
rect -313 -1793 -309 -1791
rect -303 -1793 -277 -1791
rect -269 -1793 -266 -1791
rect -247 -1793 -243 -1791
rect -237 -1793 -211 -1791
rect -203 -1793 -200 -1791
rect -158 -1794 -154 -1792
rect -148 -1794 -122 -1792
rect -114 -1794 -111 -1792
rect 27 -1803 31 -1801
rect 37 -1803 63 -1801
rect 71 -1803 74 -1801
rect 93 -1803 97 -1801
rect 103 -1803 129 -1801
rect 137 -1803 140 -1801
rect 182 -1804 186 -1802
rect 192 -1804 218 -1802
rect 226 -1804 229 -1802
rect 317 -1803 321 -1801
rect 327 -1803 353 -1801
rect 361 -1803 364 -1801
rect 396 -1802 400 -1800
rect 406 -1802 432 -1800
rect 440 -1802 443 -1800
rect 537 -1801 541 -1799
rect 547 -1801 573 -1799
rect 581 -1801 584 -1799
rect 462 -1809 466 -1807
rect 472 -1809 498 -1807
rect 506 -1809 509 -1807
rect -618 -1826 -614 -1824
rect -608 -1826 -582 -1824
rect -574 -1826 -571 -1824
rect -552 -1826 -548 -1824
rect -542 -1826 -516 -1824
rect -508 -1826 -505 -1824
rect -463 -1827 -459 -1825
rect -453 -1827 -427 -1825
rect -419 -1827 -416 -1825
rect -247 -1827 -243 -1825
rect -237 -1827 -211 -1825
rect -203 -1827 -200 -1825
rect -106 -1826 -102 -1824
rect -96 -1826 -70 -1824
rect -62 -1826 -59 -1824
rect 317 -1826 321 -1824
rect 327 -1826 353 -1824
rect 361 -1826 364 -1824
rect -181 -1834 -177 -1832
rect -171 -1834 -145 -1832
rect -137 -1834 -134 -1832
rect 93 -1837 97 -1835
rect 103 -1837 129 -1835
rect 137 -1837 140 -1835
rect 234 -1836 238 -1834
rect 244 -1836 270 -1834
rect 278 -1836 281 -1834
rect -618 -1849 -614 -1847
rect -608 -1849 -582 -1847
rect -574 -1849 -571 -1847
rect -552 -1849 -548 -1847
rect -542 -1849 -516 -1847
rect -508 -1849 -505 -1847
rect -463 -1850 -459 -1848
rect -453 -1850 -427 -1848
rect -419 -1850 -416 -1848
rect 159 -1844 163 -1842
rect 169 -1844 195 -1842
rect 203 -1844 206 -1842
rect -326 -1851 -322 -1849
rect -316 -1851 -290 -1849
rect -282 -1851 -279 -1849
rect -247 -1850 -243 -1848
rect -237 -1850 -211 -1848
rect -203 -1850 -200 -1848
rect -106 -1849 -102 -1847
rect -96 -1849 -70 -1847
rect -62 -1849 -59 -1847
rect 409 -1847 413 -1845
rect 419 -1847 445 -1845
rect 453 -1847 456 -1845
rect 507 -1852 511 -1850
rect 517 -1852 543 -1850
rect 551 -1852 554 -1850
rect -181 -1857 -177 -1855
rect -171 -1857 -145 -1855
rect -137 -1857 -134 -1855
rect 14 -1861 18 -1859
rect 24 -1861 50 -1859
rect 58 -1861 61 -1859
rect 93 -1860 97 -1858
rect 103 -1860 129 -1858
rect 137 -1860 140 -1858
rect 234 -1859 238 -1857
rect 244 -1859 270 -1857
rect 278 -1859 281 -1857
rect 159 -1867 163 -1865
rect 169 -1867 195 -1865
rect 203 -1867 206 -1865
rect 409 -1870 413 -1868
rect 419 -1870 445 -1868
rect 453 -1870 456 -1868
rect -326 -1874 -322 -1872
rect -316 -1874 -290 -1872
rect -282 -1874 -279 -1872
rect 507 -1875 511 -1873
rect 517 -1875 543 -1873
rect 551 -1875 554 -1873
rect -552 -1883 -548 -1881
rect -542 -1883 -516 -1881
rect -508 -1883 -505 -1881
rect -411 -1882 -407 -1880
rect -401 -1882 -375 -1880
rect -367 -1882 -364 -1880
rect 14 -1884 18 -1882
rect 24 -1884 50 -1882
rect 58 -1884 61 -1882
rect -486 -1890 -482 -1888
rect -476 -1890 -450 -1888
rect -442 -1890 -439 -1888
rect -234 -1895 -230 -1893
rect -224 -1895 -198 -1893
rect -190 -1895 -187 -1893
rect -136 -1900 -132 -1898
rect -126 -1900 -100 -1898
rect -92 -1900 -89 -1898
rect -631 -1907 -627 -1905
rect -621 -1907 -595 -1905
rect -587 -1907 -584 -1905
rect -552 -1906 -548 -1904
rect -542 -1906 -516 -1904
rect -508 -1906 -505 -1904
rect -411 -1905 -407 -1903
rect -401 -1905 -375 -1903
rect -367 -1905 -364 -1903
rect 106 -1905 110 -1903
rect 116 -1905 142 -1903
rect 150 -1905 153 -1903
rect 204 -1910 208 -1908
rect 214 -1910 240 -1908
rect 248 -1910 251 -1908
rect -486 -1913 -482 -1911
rect -476 -1913 -450 -1911
rect -442 -1913 -439 -1911
rect -234 -1918 -230 -1916
rect -224 -1918 -198 -1916
rect -190 -1918 -187 -1916
rect -136 -1923 -132 -1921
rect -126 -1923 -100 -1921
rect -92 -1923 -89 -1921
rect 106 -1928 110 -1926
rect 116 -1928 142 -1926
rect 150 -1928 153 -1926
rect -631 -1930 -627 -1928
rect -621 -1930 -595 -1928
rect -587 -1930 -584 -1928
rect 204 -1933 208 -1931
rect 214 -1933 240 -1931
rect 248 -1933 251 -1931
rect -539 -1951 -535 -1949
rect -529 -1951 -503 -1949
rect -495 -1951 -492 -1949
rect -441 -1956 -437 -1954
rect -431 -1956 -405 -1954
rect -397 -1956 -394 -1954
rect -539 -1974 -535 -1972
rect -529 -1974 -503 -1972
rect -495 -1974 -492 -1972
rect -441 -1979 -437 -1977
rect -431 -1979 -405 -1977
rect -397 -1979 -394 -1977
rect 451 -2039 453 -2036
rect 474 -2039 476 -2036
rect 451 -2073 453 -2047
rect 474 -2073 476 -2047
rect 525 -2069 527 -2066
rect 548 -2069 550 -2066
rect 451 -2083 453 -2079
rect 474 -2083 476 -2079
rect 259 -2093 261 -2090
rect 282 -2093 284 -2090
rect 316 -2093 318 -2090
rect 339 -2093 341 -2090
rect 396 -2091 398 -2088
rect 419 -2091 421 -2088
rect 259 -2127 261 -2101
rect 282 -2127 284 -2101
rect 316 -2127 318 -2101
rect 339 -2127 341 -2101
rect 396 -2125 398 -2099
rect 419 -2125 421 -2099
rect 525 -2103 527 -2077
rect 548 -2103 550 -2077
rect 459 -2114 461 -2111
rect 482 -2114 484 -2111
rect 525 -2113 527 -2109
rect 548 -2113 550 -2109
rect 259 -2137 261 -2133
rect 282 -2137 284 -2133
rect 316 -2137 318 -2133
rect 339 -2137 341 -2133
rect 396 -2135 398 -2131
rect 419 -2135 421 -2131
rect 459 -2148 461 -2122
rect 482 -2148 484 -2122
rect 459 -2158 461 -2154
rect 482 -2158 484 -2154
<< polycontact >>
rect -498 -471 -494 -467
rect -422 -471 -418 -467
rect -347 -471 -343 -467
rect -270 -471 -266 -467
rect -193 -471 -189 -467
rect -117 -471 -113 -467
rect -26 -471 -22 -467
rect 54 -470 58 -466
rect 133 -469 137 -465
rect 209 -468 213 -464
rect 523 -467 527 -463
rect 605 -467 609 -463
rect 685 -467 689 -463
rect 814 -468 818 -464
rect 911 -468 915 -464
rect 995 -470 999 -466
rect -504 -494 -500 -490
rect -428 -494 -424 -490
rect -353 -494 -349 -490
rect -276 -494 -272 -490
rect -199 -494 -195 -490
rect -123 -494 -119 -490
rect -32 -494 -28 -490
rect 48 -493 52 -489
rect 127 -492 131 -488
rect 203 -491 207 -487
rect 517 -490 521 -486
rect 599 -490 603 -486
rect 679 -490 683 -486
rect 808 -491 812 -487
rect 905 -491 909 -487
rect 989 -493 993 -489
rect -498 -527 -494 -523
rect -422 -527 -418 -523
rect -347 -527 -343 -523
rect -270 -527 -266 -523
rect -193 -527 -189 -523
rect -117 -527 -113 -523
rect -26 -527 -22 -523
rect 54 -526 58 -522
rect 133 -525 137 -521
rect 209 -524 213 -520
rect 523 -523 527 -519
rect 605 -523 609 -519
rect 685 -523 689 -519
rect 814 -524 818 -520
rect 911 -524 915 -520
rect 995 -526 999 -522
rect -504 -550 -500 -546
rect -428 -550 -424 -546
rect -353 -550 -349 -546
rect -276 -550 -272 -546
rect -199 -550 -195 -546
rect -123 -550 -119 -546
rect -32 -550 -28 -546
rect 48 -549 52 -545
rect 127 -548 131 -544
rect 203 -547 207 -543
rect 517 -546 521 -542
rect 599 -546 603 -542
rect 679 -546 683 -542
rect 808 -547 812 -543
rect 905 -547 909 -543
rect 989 -549 993 -545
rect 866 -649 870 -645
rect 889 -655 893 -651
rect 463 -675 467 -671
rect 61 -695 65 -691
rect 84 -701 88 -697
rect 486 -681 490 -677
rect 940 -679 944 -675
rect -388 -717 -384 -713
rect 135 -725 139 -721
rect -394 -740 -390 -736
rect -477 -745 -473 -741
rect -125 -755 -121 -751
rect -102 -749 -98 -745
rect -68 -755 -64 -751
rect -45 -749 -41 -745
rect 6 -747 10 -743
rect 29 -753 33 -749
rect 158 -731 162 -727
rect 537 -705 541 -701
rect 277 -735 281 -731
rect 300 -729 304 -725
rect 334 -735 338 -731
rect 357 -729 361 -725
rect 408 -727 412 -723
rect 431 -733 435 -729
rect 560 -711 564 -707
rect 680 -709 684 -705
rect 703 -703 707 -699
rect 737 -709 741 -705
rect 760 -703 764 -699
rect 811 -701 815 -697
rect 834 -707 838 -703
rect 963 -685 967 -681
rect 874 -724 878 -720
rect 897 -730 901 -726
rect 471 -750 475 -746
rect -483 -768 -479 -764
rect -336 -772 -332 -768
rect 69 -770 73 -766
rect -411 -780 -407 -776
rect 92 -776 96 -772
rect 494 -756 498 -752
rect -342 -795 -338 -791
rect -477 -802 -473 -798
rect -417 -803 -413 -799
rect -483 -825 -479 -821
rect -366 -846 -362 -842
rect -372 -869 -368 -865
rect -538 -928 -534 -924
rect -472 -928 -468 -924
rect -383 -929 -379 -925
rect -80 -928 -76 -924
rect -544 -951 -540 -947
rect -478 -951 -474 -947
rect -389 -952 -385 -948
rect -86 -951 -82 -947
rect 253 -947 257 -943
rect -169 -956 -165 -952
rect 247 -970 251 -966
rect -175 -979 -171 -975
rect 164 -975 168 -971
rect -472 -985 -468 -981
rect -331 -984 -327 -980
rect -28 -983 -24 -979
rect -406 -992 -402 -988
rect -103 -991 -99 -987
rect 796 -986 800 -982
rect 158 -998 162 -994
rect -551 -1009 -547 -1005
rect -478 -1008 -474 -1004
rect -337 -1007 -333 -1003
rect -34 -1006 -30 -1002
rect 305 -1002 309 -998
rect -412 -1015 -408 -1011
rect -169 -1013 -165 -1009
rect -109 -1014 -105 -1010
rect 230 -1010 234 -1006
rect 790 -1009 794 -1005
rect 707 -1014 711 -1010
rect 299 -1025 303 -1021
rect -557 -1032 -553 -1028
rect -175 -1036 -171 -1032
rect 164 -1032 168 -1028
rect 224 -1033 228 -1029
rect 701 -1037 705 -1033
rect 848 -1041 852 -1037
rect -459 -1053 -455 -1049
rect 773 -1049 777 -1045
rect -361 -1058 -357 -1054
rect -58 -1057 -54 -1053
rect 158 -1055 162 -1051
rect 842 -1064 846 -1060
rect 707 -1071 711 -1067
rect -465 -1076 -461 -1072
rect -367 -1081 -363 -1077
rect -64 -1080 -60 -1076
rect 275 -1076 279 -1072
rect 767 -1072 771 -1068
rect 701 -1094 705 -1090
rect 269 -1099 273 -1095
rect 818 -1115 822 -1111
rect -230 -1139 -226 -1135
rect -164 -1139 -160 -1135
rect -75 -1140 -71 -1136
rect 812 -1138 816 -1134
rect -236 -1162 -232 -1158
rect -170 -1162 -166 -1158
rect 103 -1158 107 -1154
rect 169 -1158 173 -1154
rect -81 -1163 -77 -1159
rect 258 -1159 262 -1155
rect 97 -1181 101 -1177
rect 163 -1181 167 -1177
rect 252 -1182 256 -1178
rect -164 -1196 -160 -1192
rect -23 -1195 -19 -1191
rect 646 -1197 650 -1193
rect 712 -1197 716 -1193
rect -98 -1203 -94 -1199
rect 801 -1198 805 -1194
rect -243 -1220 -239 -1216
rect -170 -1219 -166 -1215
rect -29 -1218 -25 -1214
rect 169 -1215 173 -1211
rect 310 -1214 314 -1210
rect -104 -1226 -100 -1222
rect 235 -1222 239 -1218
rect 640 -1220 644 -1216
rect 706 -1220 710 -1216
rect 795 -1221 799 -1217
rect -249 -1243 -245 -1239
rect 90 -1239 94 -1235
rect 163 -1238 167 -1234
rect 304 -1237 308 -1233
rect 229 -1245 233 -1241
rect 712 -1254 716 -1250
rect 853 -1253 857 -1249
rect -151 -1264 -147 -1260
rect 84 -1262 88 -1258
rect 778 -1261 782 -1257
rect -53 -1269 -49 -1265
rect 633 -1278 637 -1274
rect 706 -1277 710 -1273
rect 847 -1276 851 -1272
rect -157 -1287 -153 -1283
rect 182 -1283 186 -1279
rect -59 -1292 -55 -1288
rect 280 -1288 284 -1284
rect 772 -1284 776 -1280
rect 627 -1301 631 -1297
rect 176 -1306 180 -1302
rect 274 -1311 278 -1307
rect 725 -1322 729 -1318
rect 823 -1327 827 -1323
rect 719 -1345 723 -1341
rect 817 -1350 821 -1346
rect 499 -1509 503 -1505
rect 493 -1532 497 -1528
rect 410 -1537 414 -1533
rect -144 -1557 -140 -1553
rect 404 -1560 408 -1556
rect 196 -1567 200 -1563
rect 551 -1564 555 -1560
rect 476 -1572 480 -1568
rect -150 -1580 -146 -1576
rect -233 -1585 -229 -1581
rect 190 -1590 194 -1586
rect 545 -1587 549 -1583
rect 107 -1595 111 -1591
rect 410 -1594 414 -1590
rect 470 -1595 474 -1591
rect -239 -1608 -235 -1604
rect -449 -1613 -445 -1609
rect -92 -1612 -88 -1608
rect -167 -1620 -163 -1616
rect 101 -1618 105 -1614
rect 404 -1617 408 -1613
rect 248 -1622 252 -1618
rect 173 -1630 177 -1626
rect -455 -1636 -451 -1632
rect -98 -1635 -94 -1631
rect -538 -1641 -534 -1637
rect -233 -1642 -229 -1638
rect -173 -1643 -169 -1639
rect 521 -1638 525 -1634
rect 242 -1645 246 -1641
rect 107 -1652 111 -1648
rect 167 -1653 171 -1649
rect -544 -1664 -540 -1660
rect -397 -1668 -393 -1664
rect -239 -1665 -235 -1661
rect 515 -1661 519 -1657
rect -472 -1676 -468 -1672
rect 101 -1675 105 -1671
rect -122 -1686 -118 -1682
rect -403 -1691 -399 -1687
rect -538 -1698 -534 -1694
rect -478 -1699 -474 -1695
rect 218 -1696 222 -1692
rect -128 -1709 -124 -1705
rect -544 -1721 -540 -1717
rect 212 -1719 216 -1715
rect 349 -1720 353 -1716
rect 415 -1720 419 -1716
rect 504 -1721 508 -1717
rect -427 -1742 -423 -1738
rect 343 -1743 347 -1739
rect 409 -1743 413 -1739
rect 498 -1744 502 -1740
rect -433 -1765 -429 -1761
rect -294 -1768 -290 -1764
rect -228 -1768 -224 -1764
rect -139 -1769 -135 -1765
rect 46 -1778 50 -1774
rect 112 -1778 116 -1774
rect 201 -1779 205 -1775
rect 415 -1777 419 -1773
rect 556 -1776 560 -1772
rect 481 -1784 485 -1780
rect -300 -1791 -296 -1787
rect -234 -1791 -230 -1787
rect -145 -1792 -141 -1788
rect 40 -1801 44 -1797
rect 106 -1801 110 -1797
rect 195 -1802 199 -1798
rect 336 -1801 340 -1797
rect 409 -1800 413 -1796
rect 550 -1799 554 -1795
rect 475 -1807 479 -1803
rect -599 -1824 -595 -1820
rect -533 -1824 -529 -1820
rect -444 -1825 -440 -1821
rect -228 -1825 -224 -1821
rect -87 -1824 -83 -1820
rect 330 -1824 334 -1820
rect -162 -1832 -158 -1828
rect 112 -1835 116 -1831
rect 253 -1834 257 -1830
rect 178 -1842 182 -1838
rect -605 -1847 -601 -1843
rect -539 -1847 -535 -1843
rect -450 -1848 -446 -1844
rect -307 -1849 -303 -1845
rect -234 -1848 -230 -1844
rect -93 -1847 -89 -1843
rect 428 -1845 432 -1841
rect -168 -1855 -164 -1851
rect 526 -1850 530 -1846
rect 33 -1859 37 -1855
rect 106 -1858 110 -1854
rect 247 -1857 251 -1853
rect 172 -1865 176 -1861
rect -313 -1872 -309 -1868
rect 422 -1868 426 -1864
rect -533 -1881 -529 -1877
rect -392 -1880 -388 -1876
rect 520 -1873 524 -1869
rect 27 -1882 31 -1878
rect -467 -1888 -463 -1884
rect -215 -1893 -211 -1889
rect -612 -1905 -608 -1901
rect -539 -1904 -535 -1900
rect -398 -1903 -394 -1899
rect -117 -1898 -113 -1894
rect 125 -1903 129 -1899
rect -473 -1911 -469 -1907
rect 223 -1908 227 -1904
rect -221 -1916 -217 -1912
rect -123 -1921 -119 -1917
rect -618 -1928 -614 -1924
rect 119 -1926 123 -1922
rect 217 -1931 221 -1927
rect -520 -1949 -516 -1945
rect -422 -1954 -418 -1950
rect -526 -1972 -522 -1968
rect -428 -1977 -424 -1973
rect 447 -2064 451 -2060
rect 470 -2070 474 -2066
rect 521 -2094 525 -2090
rect 261 -2124 265 -2120
rect 284 -2118 288 -2114
rect 318 -2124 322 -2120
rect 341 -2118 345 -2114
rect 392 -2116 396 -2112
rect 415 -2122 419 -2118
rect 544 -2100 548 -2096
rect 455 -2139 459 -2135
rect 478 -2145 482 -2141
<< metal1 >>
rect 913 -144 936 -143
rect -854 -147 1001 -144
rect -854 -148 918 -147
rect -854 -149 690 -148
rect 707 -149 914 -148
rect 928 -148 1001 -147
rect 935 -149 1001 -148
rect -850 -171 844 -166
rect -850 -172 -265 -171
rect -250 -172 817 -171
rect 833 -172 844 -171
rect -839 -201 612 -194
rect -110 -202 -108 -201
rect -858 -219 53 -214
rect -858 -220 -415 -219
rect -404 -220 53 -219
rect -768 -313 130 -308
rect -768 -314 -513 -313
rect -501 -314 130 -313
rect -771 -340 685 -335
rect -771 -341 -132 -340
rect -119 -341 666 -340
rect 684 -341 685 -340
rect -769 -362 907 -359
rect -769 -363 -38 -362
rect -27 -363 907 -362
rect 567 -385 728 -384
rect 913 -385 936 -384
rect -769 -388 984 -385
rect -769 -389 37 -388
rect 49 -389 984 -388
rect 567 -390 728 -389
rect -533 -438 -527 -436
rect -457 -438 -451 -436
rect -381 -438 -376 -436
rect -306 -438 -299 -436
rect -229 -438 -222 -436
rect -152 -438 -146 -436
rect -73 -438 -55 -436
rect 18 -437 25 -435
rect 98 -436 104 -434
rect 177 -435 180 -433
rect 253 -434 494 -432
rect 253 -435 558 -434
rect 564 -435 640 -434
rect 646 -435 720 -434
rect 740 -435 852 -431
rect 177 -436 852 -435
rect 860 -436 946 -435
rect 98 -437 1411 -436
rect 18 -438 494 -437
rect -533 -439 180 -438
rect -533 -440 104 -439
rect -533 -441 25 -440
rect -533 -443 -527 -441
rect -466 -443 -451 -441
rect -390 -443 -376 -441
rect -315 -443 -299 -441
rect -238 -443 -222 -441
rect -161 -443 -146 -441
rect -85 -442 -55 -441
rect -85 -443 -78 -442
rect -73 -443 -55 -442
rect 6 -442 25 -441
rect 86 -441 104 -440
rect 165 -440 180 -439
rect 241 -439 494 -438
rect 555 -439 571 -437
rect 637 -439 656 -437
rect 717 -439 746 -437
rect 241 -440 248 -439
rect 253 -440 494 -439
rect 165 -441 172 -440
rect 177 -441 180 -440
rect 86 -442 93 -441
rect 98 -442 104 -441
rect 6 -443 13 -442
rect 18 -443 25 -442
rect -530 -444 -527 -443
rect -525 -466 -521 -465
rect -525 -470 -513 -466
rect -525 -471 -519 -470
rect -524 -501 -519 -471
rect -513 -489 -507 -478
rect -504 -490 -501 -455
rect -498 -455 -481 -451
rect -498 -467 -495 -455
rect -465 -462 -461 -443
rect -455 -444 -451 -443
rect -464 -466 -461 -462
rect -473 -470 -461 -466
rect -479 -482 -475 -478
rect -497 -486 -475 -482
rect -497 -497 -490 -486
rect -479 -489 -475 -486
rect -465 -497 -461 -470
rect -449 -466 -445 -465
rect -449 -470 -437 -466
rect -449 -471 -443 -470
rect -524 -522 -521 -501
rect -507 -502 -490 -497
rect -473 -501 -461 -497
rect -524 -526 -513 -522
rect -524 -568 -519 -526
rect -513 -545 -507 -534
rect -504 -546 -501 -502
rect -498 -523 -495 -502
rect -464 -522 -461 -501
rect -473 -526 -461 -522
rect -479 -538 -475 -534
rect -497 -542 -475 -538
rect -497 -553 -490 -542
rect -479 -545 -475 -542
rect -465 -553 -461 -526
rect -507 -558 -490 -553
rect -473 -557 -461 -553
rect -448 -501 -443 -471
rect -437 -489 -431 -478
rect -428 -490 -425 -455
rect -422 -455 -405 -451
rect -422 -467 -419 -455
rect -389 -462 -385 -443
rect -379 -444 -376 -443
rect -388 -466 -385 -462
rect -397 -470 -385 -466
rect -403 -482 -399 -478
rect -421 -486 -399 -482
rect -421 -497 -414 -486
rect -403 -489 -399 -486
rect -389 -497 -385 -470
rect -374 -466 -370 -465
rect -374 -470 -362 -466
rect -374 -471 -368 -470
rect -448 -522 -445 -501
rect -431 -502 -414 -497
rect -397 -501 -385 -497
rect -448 -526 -437 -522
rect -500 -617 -497 -558
rect -448 -568 -443 -526
rect -437 -545 -431 -534
rect -428 -546 -425 -502
rect -422 -523 -419 -502
rect -388 -522 -385 -501
rect -397 -526 -385 -522
rect -403 -538 -399 -534
rect -421 -542 -399 -538
rect -421 -553 -414 -542
rect -403 -545 -399 -542
rect -389 -553 -385 -526
rect -431 -558 -414 -553
rect -397 -557 -385 -553
rect -373 -501 -368 -471
rect -362 -489 -356 -478
rect -353 -490 -350 -455
rect -347 -455 -330 -451
rect -347 -467 -344 -455
rect -314 -462 -310 -443
rect -303 -444 -299 -443
rect -313 -466 -310 -462
rect -322 -470 -310 -466
rect -328 -482 -324 -478
rect -346 -486 -324 -482
rect -346 -497 -339 -486
rect -328 -489 -324 -486
rect -314 -497 -310 -470
rect -297 -466 -293 -465
rect -297 -470 -285 -466
rect -297 -471 -291 -470
rect -373 -522 -370 -501
rect -356 -502 -339 -497
rect -322 -501 -310 -497
rect -373 -526 -362 -522
rect -424 -590 -421 -558
rect -373 -568 -368 -526
rect -362 -545 -356 -534
rect -353 -546 -350 -502
rect -347 -523 -344 -502
rect -313 -522 -310 -501
rect -322 -526 -310 -522
rect -328 -538 -324 -534
rect -346 -542 -324 -538
rect -346 -553 -339 -542
rect -328 -545 -324 -542
rect -314 -553 -310 -526
rect -356 -558 -339 -553
rect -322 -557 -310 -553
rect -522 -621 -497 -617
rect -522 -833 -518 -621
rect -500 -625 -497 -621
rect -438 -597 -421 -590
rect -438 -642 -430 -597
rect -349 -601 -346 -558
rect -389 -606 -345 -601
rect -437 -646 -432 -642
rect -437 -662 -431 -646
rect -389 -647 -381 -606
rect -349 -608 -346 -606
rect -314 -629 -310 -557
rect -296 -501 -291 -471
rect -285 -489 -279 -478
rect -276 -490 -273 -455
rect -270 -455 -253 -451
rect -270 -467 -267 -455
rect -237 -462 -233 -443
rect -226 -444 -222 -443
rect -236 -466 -233 -462
rect -245 -470 -233 -466
rect -251 -482 -247 -478
rect -269 -486 -247 -482
rect -269 -497 -262 -486
rect -251 -489 -247 -486
rect -237 -497 -233 -470
rect -220 -466 -216 -465
rect -220 -470 -208 -466
rect -220 -471 -214 -470
rect -296 -522 -293 -501
rect -279 -502 -262 -497
rect -245 -501 -233 -497
rect -296 -526 -285 -522
rect -296 -568 -291 -526
rect -285 -545 -279 -534
rect -276 -546 -273 -502
rect -270 -523 -267 -502
rect -236 -522 -233 -501
rect -245 -526 -233 -522
rect -251 -538 -247 -534
rect -269 -542 -247 -538
rect -269 -553 -262 -542
rect -251 -545 -247 -542
rect -237 -553 -233 -526
rect -279 -558 -262 -553
rect -245 -557 -233 -553
rect -219 -501 -214 -471
rect -208 -489 -202 -478
rect -199 -490 -196 -455
rect -193 -455 -176 -451
rect -193 -467 -190 -455
rect -160 -462 -156 -443
rect -149 -444 -146 -443
rect -159 -466 -156 -462
rect -168 -470 -156 -466
rect -174 -482 -170 -478
rect -192 -486 -170 -482
rect -192 -497 -185 -486
rect -174 -489 -170 -486
rect -160 -497 -156 -470
rect -144 -466 -140 -465
rect -144 -470 -132 -466
rect -144 -471 -138 -470
rect -219 -522 -216 -501
rect -202 -502 -185 -497
rect -168 -501 -156 -497
rect -219 -526 -208 -522
rect -389 -681 -382 -647
rect -483 -685 -379 -681
rect -503 -740 -500 -693
rect -503 -744 -492 -740
rect -503 -775 -498 -744
rect -492 -763 -486 -752
rect -483 -764 -480 -685
rect -417 -694 -400 -693
rect -385 -693 -380 -685
rect -395 -694 -391 -693
rect -417 -697 -391 -694
rect -417 -713 -414 -697
rect -477 -718 -414 -713
rect -477 -741 -474 -718
rect -443 -740 -440 -724
rect -417 -734 -414 -718
rect -452 -744 -440 -740
rect -458 -756 -454 -752
rect -476 -760 -454 -756
rect -476 -771 -469 -760
rect -458 -763 -454 -760
rect -444 -771 -440 -744
rect -503 -797 -500 -775
rect -486 -776 -469 -771
rect -452 -775 -440 -771
rect -431 -775 -427 -734
rect -421 -737 -414 -734
rect -411 -716 -403 -712
rect -421 -749 -418 -737
rect -411 -740 -408 -716
rect -403 -735 -397 -724
rect -394 -736 -391 -697
rect -388 -697 -333 -693
rect -388 -713 -385 -697
rect -363 -716 -351 -712
rect -369 -728 -365 -724
rect -387 -732 -365 -728
rect -387 -743 -380 -732
rect -369 -735 -365 -732
rect -355 -743 -351 -716
rect -397 -748 -380 -743
rect -363 -747 -351 -743
rect -421 -753 -414 -749
rect -419 -755 -414 -753
rect -503 -801 -492 -797
rect -503 -832 -498 -801
rect -492 -820 -486 -809
rect -483 -821 -480 -776
rect -477 -798 -474 -776
rect -443 -797 -440 -775
rect -452 -801 -440 -797
rect -458 -813 -454 -809
rect -476 -817 -454 -813
rect -476 -828 -469 -817
rect -458 -820 -454 -817
rect -444 -828 -440 -801
rect -436 -779 -426 -775
rect -436 -823 -432 -779
rect -426 -798 -420 -787
rect -417 -799 -414 -755
rect -386 -759 -383 -748
rect -354 -756 -351 -747
rect -411 -764 -339 -759
rect -411 -776 -408 -764
rect -362 -771 -351 -767
rect -386 -779 -374 -775
rect -392 -791 -388 -787
rect -410 -795 -388 -791
rect -410 -806 -403 -795
rect -392 -798 -388 -795
rect -378 -806 -374 -779
rect -362 -802 -357 -771
rect -351 -790 -345 -779
rect -342 -791 -339 -764
rect -336 -768 -333 -697
rect -304 -767 -299 -742
rect -311 -771 -299 -767
rect -317 -783 -313 -779
rect -335 -787 -313 -783
rect -335 -798 -328 -787
rect -317 -790 -313 -787
rect -303 -798 -299 -771
rect -345 -803 -328 -798
rect -311 -802 -299 -798
rect -420 -811 -403 -806
rect -386 -810 -374 -806
rect -436 -828 -422 -823
rect -575 -839 -518 -833
rect -575 -974 -572 -839
rect -502 -842 -498 -832
rect -486 -833 -469 -828
rect -452 -832 -440 -828
rect -565 -852 -497 -842
rect -565 -923 -559 -852
rect -480 -864 -473 -833
rect -551 -871 -473 -864
rect -427 -860 -421 -828
rect -410 -830 -404 -811
rect -377 -819 -374 -810
rect -335 -823 -330 -803
rect -302 -812 -299 -802
rect -301 -819 -299 -812
rect -366 -829 -330 -823
rect -410 -836 -369 -830
rect -392 -845 -381 -841
rect -392 -860 -387 -845
rect -427 -866 -387 -860
rect -551 -910 -543 -871
rect -392 -876 -387 -866
rect -381 -864 -375 -853
rect -372 -865 -369 -836
rect -366 -842 -363 -829
rect -341 -845 -329 -841
rect -347 -857 -343 -853
rect -365 -861 -343 -857
rect -365 -872 -358 -861
rect -347 -864 -343 -861
rect -333 -861 -329 -845
rect -302 -861 -299 -819
rect -333 -866 -299 -861
rect -333 -872 -329 -866
rect -375 -877 -358 -872
rect -341 -876 -329 -872
rect -365 -880 -358 -877
rect -478 -887 -358 -880
rect -332 -885 -329 -876
rect -504 -899 -494 -890
rect -549 -915 -544 -910
rect -499 -911 -494 -899
rect -549 -918 -534 -915
rect -565 -926 -553 -923
rect -586 -979 -572 -974
rect -564 -927 -553 -926
rect -564 -958 -559 -927
rect -553 -946 -547 -935
rect -544 -947 -541 -918
rect -538 -920 -534 -918
rect -538 -924 -535 -920
rect -498 -923 -495 -911
rect -513 -927 -501 -923
rect -519 -939 -515 -935
rect -537 -943 -515 -939
rect -537 -954 -530 -943
rect -519 -946 -515 -943
rect -505 -954 -501 -927
rect -586 -1168 -581 -979
rect -564 -983 -561 -958
rect -547 -959 -530 -954
rect -513 -958 -501 -954
rect -543 -975 -539 -959
rect -505 -970 -501 -958
rect -502 -975 -501 -970
rect -498 -927 -487 -923
rect -498 -958 -493 -927
rect -487 -946 -481 -935
rect -478 -947 -475 -887
rect -472 -901 -404 -898
rect -472 -924 -469 -901
rect -412 -905 -404 -901
rect -365 -905 -358 -887
rect -438 -908 -435 -907
rect -440 -923 -435 -908
rect -412 -909 -386 -905
rect -447 -927 -435 -923
rect -412 -925 -409 -909
rect -453 -939 -449 -935
rect -471 -943 -449 -939
rect -471 -954 -464 -943
rect -453 -946 -449 -943
rect -439 -954 -435 -927
rect -577 -987 -561 -983
rect -557 -979 -539 -975
rect -577 -1004 -573 -987
rect -577 -1008 -566 -1004
rect -577 -1036 -572 -1008
rect -566 -1027 -560 -1016
rect -557 -1028 -554 -979
rect -498 -980 -495 -958
rect -481 -959 -464 -954
rect -447 -958 -435 -954
rect -551 -987 -503 -983
rect -551 -1005 -548 -987
rect -526 -1008 -514 -1004
rect -532 -1020 -528 -1016
rect -550 -1024 -528 -1020
rect -550 -1035 -543 -1024
rect -532 -1027 -528 -1024
rect -518 -1035 -514 -1008
rect -577 -1049 -570 -1036
rect -560 -1040 -543 -1035
rect -526 -1039 -514 -1035
rect -576 -1114 -570 -1049
rect -517 -1048 -514 -1039
rect -517 -1100 -513 -1048
rect -510 -1090 -503 -987
rect -498 -984 -487 -980
rect -498 -1062 -493 -984
rect -487 -1003 -481 -992
rect -478 -1004 -475 -959
rect -472 -981 -469 -959
rect -438 -980 -435 -958
rect -417 -929 -409 -925
rect -406 -928 -398 -924
rect -417 -968 -414 -929
rect -406 -959 -403 -928
rect -398 -947 -392 -936
rect -389 -948 -386 -909
rect -383 -909 -328 -905
rect -302 -909 -299 -866
rect -383 -925 -380 -909
rect -358 -928 -346 -924
rect -364 -940 -360 -936
rect -382 -944 -360 -940
rect -382 -955 -375 -944
rect -364 -947 -360 -944
rect -350 -955 -346 -928
rect -392 -960 -375 -955
rect -358 -959 -346 -955
rect -417 -971 -409 -968
rect -381 -971 -378 -960
rect -349 -968 -346 -959
rect -337 -971 -334 -964
rect -447 -984 -435 -980
rect -453 -996 -449 -992
rect -471 -1000 -449 -996
rect -471 -1011 -464 -1000
rect -453 -1003 -449 -1000
rect -439 -1011 -435 -984
rect -481 -1016 -464 -1011
rect -447 -1015 -435 -1011
rect -470 -1040 -465 -1016
rect -432 -991 -421 -987
rect -432 -1021 -427 -991
rect -421 -1010 -415 -999
rect -412 -1011 -409 -971
rect -406 -976 -334 -971
rect -406 -988 -403 -976
rect -357 -983 -346 -979
rect -381 -991 -369 -987
rect -387 -1003 -383 -999
rect -405 -1007 -383 -1003
rect -405 -1018 -398 -1007
rect -387 -1010 -383 -1007
rect -373 -1018 -369 -991
rect -357 -1014 -352 -983
rect -346 -1002 -340 -991
rect -337 -1003 -334 -976
rect -331 -980 -328 -909
rect -301 -915 -299 -909
rect -302 -950 -299 -915
rect -302 -954 -294 -950
rect -297 -979 -294 -954
rect -306 -983 -294 -979
rect -312 -995 -308 -991
rect -330 -999 -308 -995
rect -330 -1010 -323 -999
rect -312 -1002 -308 -999
rect -298 -1010 -294 -983
rect -340 -1015 -323 -1010
rect -306 -1014 -294 -1010
rect -432 -1027 -426 -1021
rect -415 -1023 -398 -1018
rect -381 -1022 -369 -1018
rect -432 -1031 -410 -1027
rect -470 -1043 -455 -1040
rect -485 -1052 -474 -1048
rect -485 -1062 -480 -1052
rect -498 -1066 -480 -1062
rect -485 -1083 -480 -1066
rect -474 -1071 -468 -1060
rect -465 -1072 -462 -1043
rect -459 -1045 -455 -1043
rect -459 -1049 -456 -1045
rect -434 -1052 -422 -1048
rect -440 -1064 -436 -1060
rect -458 -1068 -436 -1064
rect -458 -1079 -451 -1068
rect -440 -1071 -436 -1068
rect -426 -1079 -422 -1052
rect -468 -1084 -451 -1079
rect -434 -1083 -422 -1079
rect -462 -1090 -455 -1084
rect -510 -1096 -455 -1090
rect -462 -1097 -455 -1096
rect -425 -1100 -422 -1083
rect -517 -1105 -422 -1100
rect -416 -1114 -410 -1031
rect -405 -1042 -399 -1023
rect -372 -1031 -369 -1022
rect -330 -1035 -325 -1015
rect -297 -1023 -294 -1014
rect -296 -1030 -294 -1023
rect -361 -1041 -325 -1035
rect -405 -1045 -364 -1042
rect -400 -1048 -364 -1045
rect -387 -1057 -376 -1053
rect -387 -1088 -382 -1057
rect -376 -1076 -370 -1065
rect -367 -1077 -364 -1048
rect -361 -1054 -358 -1041
rect -297 -1053 -294 -1030
rect -336 -1057 -294 -1053
rect -328 -1058 -294 -1057
rect -342 -1069 -338 -1065
rect -360 -1073 -338 -1069
rect -360 -1084 -353 -1073
rect -342 -1076 -338 -1073
rect -328 -1084 -324 -1058
rect -387 -1114 -381 -1088
rect -370 -1089 -353 -1084
rect -336 -1088 -324 -1084
rect -576 -1121 -381 -1114
rect -576 -1123 -573 -1121
rect -561 -1122 -381 -1121
rect -561 -1123 -382 -1122
rect -537 -1137 -380 -1129
rect -586 -1174 -493 -1168
rect -498 -1547 -493 -1174
rect -388 -1500 -380 -1137
rect -367 -1179 -361 -1089
rect -327 -1097 -324 -1088
rect -272 -1179 -269 -558
rect -219 -568 -214 -526
rect -208 -545 -202 -534
rect -199 -546 -196 -502
rect -193 -523 -190 -502
rect -159 -522 -156 -501
rect -168 -526 -156 -522
rect -174 -538 -170 -534
rect -192 -542 -170 -538
rect -192 -553 -185 -542
rect -174 -545 -170 -542
rect -160 -553 -156 -526
rect -202 -558 -185 -553
rect -168 -557 -156 -553
rect -143 -501 -138 -471
rect -132 -489 -126 -478
rect -123 -490 -120 -455
rect -117 -455 -100 -451
rect -117 -467 -114 -455
rect -84 -462 -80 -443
rect -83 -466 -80 -462
rect -92 -470 -80 -466
rect -98 -482 -94 -478
rect -116 -486 -94 -482
rect -116 -497 -109 -486
rect -98 -489 -94 -486
rect -84 -497 -80 -470
rect -143 -522 -140 -501
rect -126 -502 -109 -497
rect -92 -501 -80 -497
rect -143 -526 -132 -522
rect -195 -594 -192 -558
rect -143 -568 -138 -526
rect -132 -545 -126 -534
rect -123 -546 -120 -502
rect -117 -523 -114 -502
rect -83 -522 -80 -501
rect -92 -526 -80 -522
rect -98 -538 -94 -534
rect -116 -542 -94 -538
rect -116 -553 -109 -542
rect -98 -545 -94 -542
rect -84 -553 -80 -526
rect -126 -558 -109 -553
rect -92 -557 -80 -553
rect -196 -845 -192 -594
rect -119 -685 -116 -558
rect -73 -655 -67 -443
rect -58 -444 -55 -443
rect -53 -466 -49 -465
rect -53 -470 -41 -466
rect -53 -471 -47 -470
rect -52 -501 -47 -471
rect -41 -489 -35 -478
rect -32 -490 -29 -455
rect -26 -455 -9 -451
rect -26 -467 -23 -455
rect 7 -466 11 -443
rect -1 -470 11 -466
rect 27 -465 31 -464
rect 27 -469 39 -465
rect 27 -470 33 -469
rect -7 -482 -3 -478
rect -25 -486 -3 -482
rect -25 -497 -18 -486
rect -7 -489 -3 -486
rect 7 -497 11 -470
rect -52 -522 -49 -501
rect -35 -502 -18 -497
rect -1 -501 11 -497
rect -52 -526 -41 -522
rect -52 -568 -47 -526
rect -41 -545 -35 -534
rect -32 -546 -29 -502
rect -26 -523 -23 -502
rect 8 -522 11 -501
rect -1 -526 11 -522
rect -7 -538 -3 -534
rect -25 -542 -3 -538
rect -25 -553 -18 -542
rect -7 -545 -3 -542
rect 7 -553 11 -526
rect -35 -558 -18 -553
rect -1 -557 11 -553
rect 28 -500 33 -470
rect 39 -488 45 -477
rect 48 -489 51 -454
rect 54 -454 71 -450
rect 54 -466 57 -454
rect 87 -461 91 -442
rect 88 -465 91 -461
rect 79 -469 91 -465
rect 106 -464 110 -463
rect 106 -468 118 -464
rect 106 -469 112 -468
rect 73 -481 77 -477
rect 55 -485 77 -481
rect 55 -496 62 -485
rect 73 -488 77 -485
rect 87 -496 91 -469
rect 28 -521 31 -500
rect 45 -501 62 -496
rect 79 -500 91 -496
rect 28 -525 39 -521
rect -28 -654 -25 -558
rect 28 -567 33 -525
rect 39 -544 45 -533
rect 48 -545 51 -501
rect 54 -522 57 -501
rect 88 -521 91 -500
rect 79 -525 91 -521
rect 73 -537 77 -533
rect 55 -541 77 -537
rect 55 -552 62 -541
rect 73 -544 77 -541
rect 87 -552 91 -525
rect 45 -557 62 -552
rect 79 -556 91 -552
rect 107 -499 112 -469
rect 118 -487 124 -476
rect 127 -488 130 -453
rect 133 -453 150 -449
rect 133 -465 136 -453
rect 166 -460 170 -441
rect 167 -464 170 -460
rect 158 -468 170 -464
rect 182 -463 186 -462
rect 182 -467 194 -463
rect 182 -468 188 -467
rect 152 -480 156 -476
rect 134 -484 156 -480
rect 134 -495 141 -484
rect 152 -487 156 -484
rect 166 -495 170 -468
rect 107 -520 110 -499
rect 124 -500 141 -495
rect 158 -499 170 -495
rect 107 -524 118 -520
rect 52 -615 55 -557
rect 107 -566 112 -524
rect 118 -543 124 -532
rect 127 -544 130 -500
rect 133 -521 136 -500
rect 167 -520 170 -499
rect 158 -524 170 -520
rect 152 -536 156 -532
rect 134 -540 156 -536
rect 134 -551 141 -540
rect 152 -543 156 -540
rect 166 -551 170 -524
rect 124 -556 141 -551
rect 158 -555 170 -551
rect 183 -498 188 -468
rect 194 -486 200 -475
rect 203 -487 206 -452
rect 209 -452 226 -448
rect 209 -464 212 -452
rect 242 -459 246 -440
rect 243 -463 246 -459
rect 234 -467 246 -463
rect 228 -479 232 -475
rect 210 -483 232 -479
rect 210 -494 217 -483
rect 228 -486 232 -483
rect 242 -494 246 -467
rect 183 -519 186 -498
rect 200 -499 217 -494
rect 234 -498 246 -494
rect 183 -523 194 -519
rect 131 -606 134 -556
rect 183 -565 188 -523
rect 194 -542 200 -531
rect 203 -543 206 -499
rect 209 -520 212 -499
rect 243 -519 246 -498
rect 234 -523 246 -519
rect 228 -535 232 -531
rect 210 -539 232 -535
rect 210 -550 217 -539
rect 228 -542 232 -539
rect 242 -550 246 -523
rect 200 -555 217 -550
rect 234 -554 246 -550
rect -12 -618 55 -615
rect -12 -654 -9 -618
rect 207 -610 210 -555
rect 254 -595 260 -440
rect 496 -462 500 -461
rect 496 -466 508 -462
rect 496 -467 502 -466
rect 497 -497 502 -467
rect 508 -485 514 -474
rect 517 -486 520 -451
rect 523 -451 540 -447
rect 523 -463 526 -451
rect 556 -458 560 -439
rect 557 -462 560 -458
rect 548 -466 560 -462
rect 542 -478 546 -474
rect 524 -482 546 -478
rect 524 -493 531 -482
rect 542 -485 546 -482
rect 556 -493 560 -466
rect 578 -462 582 -461
rect 578 -466 590 -462
rect 578 -467 584 -466
rect 497 -518 500 -497
rect 514 -498 531 -493
rect 548 -497 560 -493
rect 497 -522 508 -518
rect 497 -564 502 -522
rect 508 -541 514 -530
rect 517 -542 520 -498
rect 523 -519 526 -498
rect 557 -518 560 -497
rect 548 -522 560 -518
rect 542 -534 546 -530
rect 524 -538 546 -534
rect 524 -549 531 -538
rect 542 -541 546 -538
rect 556 -549 560 -522
rect 514 -554 531 -549
rect 548 -553 560 -549
rect 579 -497 584 -467
rect 590 -485 596 -474
rect 599 -486 602 -451
rect 605 -451 622 -447
rect 605 -463 608 -451
rect 638 -458 642 -439
rect 639 -462 642 -458
rect 630 -466 642 -462
rect 624 -478 628 -474
rect 606 -482 628 -478
rect 606 -493 613 -482
rect 624 -485 628 -482
rect 638 -493 642 -466
rect 658 -462 662 -461
rect 658 -466 670 -462
rect 658 -467 664 -466
rect 579 -518 582 -497
rect 596 -498 613 -493
rect 630 -497 642 -493
rect 579 -522 590 -518
rect 254 -603 476 -595
rect 470 -608 476 -603
rect 337 -610 476 -608
rect 521 -601 524 -554
rect 579 -564 584 -522
rect 590 -541 596 -530
rect 599 -542 602 -498
rect 605 -519 608 -498
rect 639 -518 642 -497
rect 630 -522 642 -518
rect 624 -534 628 -530
rect 606 -538 628 -534
rect 606 -549 613 -538
rect 624 -541 628 -538
rect 638 -549 642 -522
rect 596 -554 613 -549
rect 630 -553 642 -549
rect 659 -497 664 -467
rect 670 -485 676 -474
rect 679 -486 682 -451
rect 685 -451 702 -447
rect 685 -463 688 -451
rect 718 -458 722 -439
rect 719 -462 722 -458
rect 710 -466 722 -462
rect 704 -478 708 -474
rect 686 -482 708 -478
rect 686 -493 693 -482
rect 704 -485 708 -482
rect 718 -493 722 -466
rect 659 -518 662 -497
rect 676 -498 693 -493
rect 710 -497 722 -493
rect 659 -522 670 -518
rect -72 -663 -59 -655
rect -28 -657 -21 -654
rect -65 -669 -59 -663
rect -156 -686 -116 -685
rect -165 -691 -116 -686
rect -165 -692 -125 -691
rect -165 -804 -162 -692
rect -26 -699 -21 -657
rect -147 -705 -21 -699
rect -14 -692 -8 -654
rect 60 -661 104 -658
rect 60 -662 95 -661
rect 60 -670 64 -662
rect 91 -670 95 -662
rect 72 -676 83 -672
rect 76 -687 80 -676
rect 76 -689 96 -687
rect -14 -695 61 -692
rect 76 -694 122 -689
rect -147 -778 -141 -705
rect -132 -714 -65 -712
rect -59 -714 -24 -712
rect -132 -715 -24 -714
rect -132 -716 -97 -715
rect -132 -724 -128 -716
rect -101 -724 -97 -716
rect -120 -730 -109 -726
rect -117 -741 -113 -730
rect -75 -716 -40 -715
rect -75 -724 -71 -716
rect -44 -724 -40 -716
rect -63 -730 -52 -726
rect -60 -741 -56 -730
rect -133 -746 -113 -741
rect -132 -748 -113 -746
rect -132 -752 -128 -748
rect -76 -746 -56 -741
rect -14 -743 -10 -695
rect 52 -701 84 -698
rect 5 -713 49 -710
rect 5 -714 40 -713
rect 5 -722 9 -714
rect 36 -722 40 -714
rect 17 -728 28 -724
rect 21 -739 25 -728
rect 21 -742 41 -739
rect 52 -742 57 -701
rect 91 -704 96 -694
rect 72 -710 83 -704
rect 60 -716 64 -710
rect 60 -721 95 -716
rect 116 -722 122 -694
rect 134 -691 178 -688
rect 134 -692 169 -691
rect 134 -700 138 -692
rect 165 -700 169 -692
rect 146 -706 157 -702
rect 150 -717 154 -706
rect 116 -725 135 -722
rect 150 -724 170 -717
rect 123 -731 158 -728
rect -33 -744 -10 -743
rect -98 -748 -56 -746
rect -98 -749 -71 -748
rect -33 -746 6 -744
rect -41 -747 6 -746
rect 21 -745 57 -742
rect 21 -746 41 -745
rect -41 -749 -30 -747
rect -133 -758 -128 -752
rect -76 -752 -71 -749
rect -121 -755 -71 -752
rect -14 -752 29 -750
rect -64 -753 29 -752
rect -64 -755 -10 -753
rect -76 -758 -71 -755
rect -120 -764 -109 -758
rect -63 -764 -52 -758
rect -101 -770 -97 -764
rect -44 -770 -40 -764
rect -132 -772 -97 -770
rect -75 -772 -40 -770
rect -132 -775 -24 -772
rect -14 -773 -10 -755
rect 36 -756 41 -746
rect 17 -762 28 -756
rect 5 -767 9 -762
rect 5 -770 39 -767
rect 52 -767 57 -745
rect 68 -736 112 -733
rect 68 -737 103 -736
rect 68 -745 72 -737
rect 99 -745 103 -737
rect 80 -751 91 -747
rect 84 -762 88 -751
rect 84 -763 104 -762
rect 123 -763 129 -731
rect 165 -734 170 -724
rect 52 -770 69 -767
rect 84 -769 129 -763
rect 146 -740 157 -734
rect 134 -746 138 -740
rect 134 -751 169 -746
rect -14 -776 92 -773
rect -14 -778 -8 -776
rect -147 -783 -8 -778
rect 99 -779 104 -769
rect 80 -785 91 -779
rect 68 -791 72 -785
rect 134 -790 140 -751
rect 102 -791 140 -790
rect 68 -796 140 -791
rect -165 -809 -123 -804
rect -129 -838 -123 -809
rect -92 -827 -86 -806
rect 109 -809 122 -802
rect -92 -833 -74 -827
rect -130 -841 -86 -838
rect -197 -853 -192 -845
rect -197 -858 -121 -853
rect -130 -867 -122 -858
rect -92 -863 -86 -841
rect -129 -873 -123 -867
rect -92 -871 -87 -863
rect -81 -892 -74 -833
rect 110 -869 118 -809
rect 206 -855 211 -610
rect 337 -614 475 -610
rect 337 -649 343 -614
rect 521 -617 525 -601
rect 603 -605 606 -554
rect 659 -564 664 -522
rect 670 -541 676 -530
rect 679 -542 682 -498
rect 685 -519 688 -498
rect 719 -518 722 -497
rect 710 -522 722 -518
rect 704 -534 708 -530
rect 686 -538 708 -534
rect 686 -549 693 -538
rect 704 -541 708 -538
rect 718 -549 722 -522
rect 676 -554 693 -549
rect 710 -553 722 -549
rect 397 -618 527 -617
rect 376 -622 527 -618
rect 376 -679 381 -622
rect 602 -625 606 -605
rect 683 -625 686 -554
rect 489 -626 606 -625
rect 394 -627 606 -626
rect 255 -685 381 -679
rect 388 -630 606 -627
rect 636 -628 686 -625
rect 740 -623 746 -439
rect 846 -438 1411 -437
rect 846 -440 863 -438
rect 943 -439 1411 -438
rect 943 -440 971 -439
rect 1022 -440 1411 -439
rect 787 -463 791 -462
rect 787 -467 799 -463
rect 787 -468 793 -467
rect 788 -498 793 -468
rect 799 -486 805 -475
rect 808 -487 811 -452
rect 814 -452 831 -448
rect 814 -464 817 -452
rect 847 -459 851 -440
rect 848 -463 851 -459
rect 839 -467 851 -463
rect 833 -479 837 -475
rect 815 -483 837 -479
rect 815 -494 822 -483
rect 833 -486 837 -483
rect 847 -494 851 -467
rect 884 -463 888 -462
rect 884 -467 896 -463
rect 884 -468 890 -467
rect 788 -519 791 -498
rect 805 -499 822 -494
rect 839 -498 851 -494
rect 788 -523 799 -519
rect 788 -565 793 -523
rect 799 -542 805 -531
rect 808 -543 811 -499
rect 814 -520 817 -499
rect 848 -519 851 -498
rect 839 -523 851 -519
rect 833 -535 837 -531
rect 815 -539 837 -535
rect 815 -550 822 -539
rect 833 -542 837 -539
rect 847 -550 851 -523
rect 805 -555 822 -550
rect 839 -554 851 -550
rect 885 -498 890 -468
rect 896 -486 902 -475
rect 905 -487 908 -452
rect 911 -452 928 -448
rect 911 -464 914 -452
rect 944 -459 948 -440
rect 1024 -441 1411 -440
rect 945 -463 948 -459
rect 936 -467 948 -463
rect 930 -479 934 -475
rect 912 -483 934 -479
rect 912 -494 919 -483
rect 930 -486 934 -483
rect 944 -494 948 -467
rect 968 -465 972 -464
rect 968 -469 980 -465
rect 968 -470 974 -469
rect 885 -519 888 -498
rect 902 -499 919 -494
rect 936 -498 948 -494
rect 885 -523 896 -519
rect 812 -592 815 -555
rect 885 -565 890 -523
rect 896 -542 902 -531
rect 905 -543 908 -499
rect 911 -520 914 -499
rect 945 -519 948 -498
rect 936 -523 948 -519
rect 930 -535 934 -531
rect 912 -539 934 -535
rect 912 -550 919 -539
rect 930 -542 934 -539
rect 944 -550 948 -523
rect 902 -555 919 -550
rect 936 -554 948 -550
rect 969 -500 974 -470
rect 980 -488 986 -477
rect 989 -489 992 -452
rect 995 -454 1006 -450
rect 995 -466 998 -454
rect 1028 -461 1032 -441
rect 1029 -465 1032 -461
rect 1020 -469 1032 -465
rect 1014 -481 1018 -477
rect 996 -485 1018 -481
rect 996 -496 1003 -485
rect 1014 -488 1018 -485
rect 1028 -496 1032 -469
rect 969 -521 972 -500
rect 986 -501 1003 -496
rect 1020 -500 1032 -496
rect 969 -525 980 -521
rect 388 -672 394 -630
rect 462 -641 506 -638
rect 462 -642 497 -641
rect 462 -650 466 -642
rect 493 -650 497 -642
rect 474 -656 485 -652
rect 478 -667 482 -656
rect 478 -669 498 -667
rect 388 -675 463 -672
rect 478 -674 524 -669
rect 255 -758 261 -685
rect 270 -694 337 -692
rect 343 -694 378 -692
rect 270 -695 378 -694
rect 270 -696 305 -695
rect 270 -704 274 -696
rect 301 -704 305 -696
rect 282 -710 293 -706
rect 285 -721 289 -710
rect 327 -696 362 -695
rect 327 -704 331 -696
rect 358 -704 362 -696
rect 339 -710 350 -706
rect 342 -721 346 -710
rect 269 -726 289 -721
rect 270 -728 289 -726
rect 270 -732 274 -728
rect 326 -726 346 -721
rect 388 -723 392 -675
rect 454 -681 486 -678
rect 407 -693 451 -690
rect 407 -694 442 -693
rect 407 -702 411 -694
rect 438 -702 442 -694
rect 419 -708 430 -704
rect 423 -719 427 -708
rect 423 -722 443 -719
rect 454 -722 459 -681
rect 493 -684 498 -674
rect 474 -690 485 -684
rect 462 -696 466 -690
rect 462 -701 497 -696
rect 518 -702 524 -674
rect 536 -671 580 -668
rect 536 -672 571 -671
rect 536 -680 540 -672
rect 567 -680 571 -672
rect 548 -686 559 -682
rect 552 -697 556 -686
rect 518 -705 537 -702
rect 552 -704 572 -697
rect 525 -711 560 -708
rect 369 -724 392 -723
rect 304 -728 346 -726
rect 304 -729 331 -728
rect 369 -726 408 -724
rect 361 -727 408 -726
rect 423 -725 459 -722
rect 423 -726 443 -725
rect 361 -729 372 -727
rect 269 -738 274 -732
rect 326 -732 331 -729
rect 281 -735 331 -732
rect 388 -732 431 -730
rect 338 -733 431 -732
rect 338 -735 392 -733
rect 326 -738 331 -735
rect 282 -744 293 -738
rect 339 -744 350 -738
rect 301 -750 305 -744
rect 358 -750 362 -744
rect 270 -752 305 -750
rect 327 -752 362 -750
rect 270 -755 378 -752
rect 388 -753 392 -735
rect 438 -736 443 -726
rect 419 -742 430 -736
rect 407 -747 411 -742
rect 407 -750 441 -747
rect 454 -747 459 -725
rect 470 -716 514 -713
rect 470 -717 505 -716
rect 470 -725 474 -717
rect 501 -725 505 -717
rect 482 -731 493 -727
rect 486 -742 490 -731
rect 486 -743 506 -742
rect 525 -743 531 -711
rect 567 -714 572 -704
rect 454 -750 471 -747
rect 486 -749 531 -743
rect 548 -720 559 -714
rect 536 -726 540 -720
rect 536 -731 571 -726
rect 388 -756 494 -753
rect 388 -758 394 -756
rect 255 -763 394 -758
rect 501 -759 506 -749
rect 482 -765 493 -759
rect 470 -771 474 -765
rect 536 -770 542 -731
rect 504 -771 542 -770
rect 470 -776 542 -771
rect 206 -859 246 -855
rect 310 -856 316 -786
rect 206 -860 211 -859
rect 110 -874 210 -869
rect 204 -892 210 -874
rect -175 -896 -71 -892
rect -195 -951 -192 -904
rect -195 -955 -184 -951
rect -195 -986 -190 -955
rect -184 -974 -178 -963
rect -175 -975 -172 -896
rect -109 -905 -92 -904
rect -77 -904 -72 -896
rect 241 -890 246 -859
rect 249 -865 316 -856
rect 514 -789 524 -782
rect 252 -870 259 -865
rect 514 -867 517 -789
rect 636 -847 639 -628
rect 779 -596 815 -592
rect 779 -653 784 -596
rect 812 -597 815 -596
rect 909 -600 912 -555
rect 969 -567 974 -525
rect 980 -544 986 -533
rect 989 -545 992 -501
rect 995 -522 998 -501
rect 1029 -521 1032 -500
rect 1020 -525 1032 -521
rect 1014 -537 1018 -533
rect 996 -541 1018 -537
rect 996 -552 1003 -541
rect 1014 -544 1018 -541
rect 1028 -552 1032 -525
rect 986 -557 1003 -552
rect 1020 -556 1032 -552
rect 797 -601 912 -600
rect 658 -659 784 -653
rect 791 -604 912 -601
rect 791 -646 797 -604
rect 865 -615 909 -612
rect 865 -616 900 -615
rect 865 -624 869 -616
rect 896 -624 900 -616
rect 877 -630 888 -626
rect 881 -641 885 -630
rect 881 -643 901 -641
rect 791 -649 866 -646
rect 881 -648 927 -643
rect 658 -732 664 -659
rect 673 -668 740 -666
rect 746 -668 781 -666
rect 673 -669 781 -668
rect 673 -670 708 -669
rect 673 -678 677 -670
rect 704 -678 708 -670
rect 685 -684 696 -680
rect 688 -695 692 -684
rect 730 -670 765 -669
rect 730 -678 734 -670
rect 761 -678 765 -670
rect 742 -684 753 -680
rect 745 -695 749 -684
rect 672 -700 692 -695
rect 673 -702 692 -700
rect 673 -706 677 -702
rect 729 -700 749 -695
rect 791 -697 795 -649
rect 857 -655 889 -652
rect 810 -667 854 -664
rect 810 -668 845 -667
rect 810 -676 814 -668
rect 841 -676 845 -668
rect 822 -682 833 -678
rect 826 -693 830 -682
rect 826 -696 846 -693
rect 857 -696 862 -655
rect 896 -658 901 -648
rect 877 -664 888 -658
rect 865 -670 869 -664
rect 865 -675 900 -670
rect 921 -676 927 -648
rect 939 -645 983 -642
rect 939 -646 974 -645
rect 939 -654 943 -646
rect 970 -654 974 -646
rect 951 -660 962 -656
rect 955 -671 959 -660
rect 921 -679 940 -676
rect 955 -678 975 -671
rect 928 -685 963 -682
rect 772 -698 795 -697
rect 707 -702 749 -700
rect 707 -703 734 -702
rect 772 -700 811 -698
rect 764 -701 811 -700
rect 826 -699 862 -696
rect 826 -700 846 -699
rect 764 -703 775 -701
rect 672 -712 677 -706
rect 729 -706 734 -703
rect 684 -709 734 -706
rect 791 -706 834 -704
rect 741 -707 834 -706
rect 741 -709 795 -707
rect 729 -712 734 -709
rect 685 -718 696 -712
rect 742 -718 753 -712
rect 704 -724 708 -718
rect 761 -724 765 -718
rect 673 -726 708 -724
rect 730 -726 765 -724
rect 673 -729 781 -726
rect 791 -727 795 -709
rect 841 -710 846 -700
rect 822 -716 833 -710
rect 810 -721 814 -716
rect 810 -724 844 -721
rect 857 -721 862 -699
rect 873 -690 917 -687
rect 873 -691 908 -690
rect 873 -699 877 -691
rect 904 -699 908 -691
rect 885 -705 896 -701
rect 889 -716 893 -705
rect 889 -717 909 -716
rect 928 -717 934 -685
rect 970 -688 975 -678
rect 857 -724 874 -721
rect 889 -723 934 -717
rect 951 -694 962 -688
rect 939 -700 943 -694
rect 939 -705 974 -700
rect 791 -730 897 -727
rect 791 -732 797 -730
rect 658 -737 797 -732
rect 904 -733 909 -723
rect 885 -739 896 -733
rect 873 -745 877 -739
rect 939 -744 945 -705
rect 907 -745 945 -744
rect 873 -750 945 -745
rect 713 -828 719 -760
rect 917 -763 927 -756
rect 713 -835 814 -828
rect 636 -850 792 -847
rect 636 -851 639 -850
rect 252 -877 260 -870
rect 514 -873 755 -867
rect -87 -905 -83 -904
rect -109 -908 -83 -905
rect -109 -924 -106 -908
rect -169 -929 -106 -924
rect -169 -952 -166 -929
rect -135 -951 -132 -935
rect -109 -945 -106 -929
rect -144 -955 -132 -951
rect -150 -967 -146 -963
rect -168 -971 -146 -967
rect -168 -982 -161 -971
rect -150 -974 -146 -971
rect -136 -982 -132 -955
rect -195 -1008 -192 -986
rect -178 -987 -161 -982
rect -144 -986 -132 -982
rect -123 -986 -119 -945
rect -113 -948 -106 -945
rect -103 -927 -95 -923
rect -113 -960 -110 -948
rect -103 -951 -100 -927
rect -95 -946 -89 -935
rect -86 -947 -83 -908
rect -80 -908 -25 -904
rect -80 -924 -77 -908
rect -55 -927 -43 -923
rect -61 -939 -57 -935
rect -79 -943 -57 -939
rect -79 -954 -72 -943
rect -61 -946 -57 -943
rect -47 -954 -43 -927
rect -89 -959 -72 -954
rect -55 -958 -43 -954
rect -113 -964 -106 -960
rect -111 -966 -106 -964
rect -195 -1012 -184 -1008
rect -195 -1043 -190 -1012
rect -184 -1031 -178 -1020
rect -175 -1032 -172 -987
rect -169 -1009 -166 -987
rect -135 -1008 -132 -986
rect -144 -1012 -132 -1008
rect -150 -1024 -146 -1020
rect -168 -1028 -146 -1024
rect -168 -1039 -161 -1028
rect -150 -1031 -146 -1028
rect -136 -1039 -132 -1012
rect -128 -990 -118 -986
rect -128 -1034 -124 -990
rect -118 -1009 -112 -998
rect -109 -1010 -106 -966
rect -78 -970 -75 -959
rect -46 -967 -43 -958
rect -103 -975 -31 -970
rect -103 -987 -100 -975
rect -54 -982 -43 -978
rect -78 -990 -66 -986
rect -84 -1002 -80 -998
rect -102 -1006 -80 -1002
rect -102 -1017 -95 -1006
rect -84 -1009 -80 -1006
rect -70 -1017 -66 -990
rect -54 -1013 -49 -982
rect -43 -1001 -37 -990
rect -34 -1002 -31 -975
rect -28 -979 -25 -908
rect 252 -911 259 -877
rect 158 -915 262 -911
rect 747 -915 752 -873
rect 4 -978 9 -953
rect -3 -982 9 -978
rect -9 -994 -5 -990
rect -27 -998 -5 -994
rect -27 -1009 -20 -998
rect -9 -1001 -5 -998
rect 5 -1009 9 -982
rect -37 -1014 -20 -1009
rect -3 -1013 9 -1009
rect -112 -1022 -95 -1017
rect -78 -1021 -66 -1017
rect -128 -1039 -114 -1034
rect -194 -1053 -190 -1043
rect -178 -1044 -161 -1039
rect -144 -1043 -132 -1039
rect -257 -1063 -189 -1053
rect -257 -1134 -251 -1063
rect -172 -1075 -165 -1044
rect -243 -1082 -165 -1075
rect -119 -1071 -113 -1039
rect -102 -1041 -96 -1022
rect -69 -1030 -66 -1021
rect -27 -1034 -22 -1014
rect 6 -1023 9 -1013
rect 7 -1030 9 -1023
rect -58 -1040 -22 -1034
rect -102 -1047 -61 -1041
rect -84 -1056 -73 -1052
rect -84 -1071 -79 -1056
rect -119 -1077 -79 -1071
rect -243 -1121 -235 -1082
rect -84 -1087 -79 -1077
rect -73 -1075 -67 -1064
rect -64 -1076 -61 -1047
rect -58 -1053 -55 -1040
rect -33 -1056 -21 -1052
rect -39 -1068 -35 -1064
rect -57 -1072 -35 -1068
rect -57 -1083 -50 -1072
rect -39 -1075 -35 -1072
rect -25 -1072 -21 -1056
rect 6 -1072 9 -1030
rect 138 -970 141 -923
rect 138 -974 149 -970
rect 138 -1005 143 -974
rect 149 -993 155 -982
rect 158 -994 161 -915
rect 224 -924 241 -923
rect 256 -923 261 -915
rect 246 -924 250 -923
rect 224 -927 250 -924
rect 224 -943 227 -927
rect 164 -948 227 -943
rect 164 -971 167 -948
rect 198 -970 201 -954
rect 224 -964 227 -948
rect 189 -974 201 -970
rect 183 -986 187 -982
rect 165 -990 187 -986
rect 165 -1001 172 -990
rect 183 -993 187 -990
rect 197 -1001 201 -974
rect 138 -1027 141 -1005
rect 155 -1006 172 -1001
rect 189 -1005 201 -1001
rect 210 -1005 214 -964
rect 220 -967 227 -964
rect 230 -946 238 -942
rect 220 -979 223 -967
rect 230 -970 233 -946
rect 238 -965 244 -954
rect 247 -966 250 -927
rect 253 -927 308 -923
rect 253 -943 256 -927
rect 278 -946 290 -942
rect 272 -958 276 -954
rect 254 -962 276 -958
rect 254 -973 261 -962
rect 272 -965 276 -962
rect 286 -973 290 -946
rect 244 -978 261 -973
rect 278 -977 290 -973
rect 220 -983 227 -979
rect 222 -985 227 -983
rect 138 -1031 149 -1027
rect 138 -1062 143 -1031
rect 149 -1050 155 -1039
rect 158 -1051 161 -1006
rect 164 -1028 167 -1006
rect 198 -1027 201 -1005
rect 189 -1031 201 -1027
rect 183 -1043 187 -1039
rect 165 -1047 187 -1043
rect 165 -1058 172 -1047
rect 183 -1050 187 -1047
rect 197 -1058 201 -1031
rect 205 -1009 215 -1005
rect 205 -1053 209 -1009
rect 215 -1028 221 -1017
rect 224 -1029 227 -985
rect 255 -989 258 -978
rect 287 -986 290 -977
rect 230 -994 302 -989
rect 230 -1006 233 -994
rect 279 -1001 290 -997
rect 255 -1009 267 -1005
rect 249 -1021 253 -1017
rect 231 -1025 253 -1021
rect 231 -1036 238 -1025
rect 249 -1028 253 -1025
rect 263 -1036 267 -1009
rect 279 -1032 284 -1001
rect 290 -1020 296 -1009
rect 299 -1021 302 -994
rect 305 -998 308 -927
rect 747 -931 753 -915
rect 784 -929 789 -850
rect 795 -916 803 -835
rect 795 -950 802 -916
rect 701 -954 805 -950
rect 337 -997 342 -972
rect 330 -1001 342 -997
rect 324 -1013 328 -1009
rect 306 -1017 328 -1013
rect 306 -1028 313 -1017
rect 324 -1020 328 -1017
rect 338 -1028 342 -1001
rect 296 -1033 313 -1028
rect 330 -1032 342 -1028
rect 221 -1041 238 -1036
rect 255 -1040 267 -1036
rect 205 -1058 219 -1053
rect 139 -1072 143 -1062
rect 155 -1063 172 -1058
rect 189 -1062 201 -1058
rect -25 -1077 9 -1072
rect -25 -1083 -21 -1077
rect -67 -1088 -50 -1083
rect -33 -1087 -21 -1083
rect -57 -1091 -50 -1088
rect -170 -1098 -50 -1091
rect -24 -1096 -21 -1087
rect -196 -1110 -186 -1101
rect -241 -1126 -236 -1121
rect -191 -1122 -186 -1110
rect -241 -1129 -226 -1126
rect -257 -1137 -245 -1134
rect -369 -1211 -361 -1179
rect -280 -1185 -269 -1179
rect -256 -1138 -245 -1137
rect -256 -1169 -251 -1138
rect -245 -1157 -239 -1146
rect -236 -1158 -233 -1129
rect -230 -1131 -226 -1129
rect -230 -1135 -227 -1131
rect -190 -1134 -187 -1122
rect -205 -1138 -193 -1134
rect -211 -1150 -207 -1146
rect -229 -1154 -207 -1150
rect -229 -1165 -222 -1154
rect -211 -1157 -207 -1154
rect -197 -1165 -193 -1138
rect -369 -1409 -362 -1211
rect -371 -1418 -362 -1409
rect -371 -1426 -363 -1418
rect -280 -1425 -276 -1185
rect -256 -1194 -253 -1169
rect -239 -1170 -222 -1165
rect -205 -1169 -193 -1165
rect -235 -1186 -231 -1170
rect -197 -1181 -193 -1169
rect -194 -1186 -193 -1181
rect -190 -1138 -179 -1134
rect -190 -1169 -185 -1138
rect -179 -1157 -173 -1146
rect -170 -1158 -167 -1098
rect -164 -1112 -96 -1109
rect -164 -1135 -161 -1112
rect -104 -1116 -96 -1112
rect -57 -1116 -50 -1098
rect -130 -1119 -127 -1118
rect -132 -1134 -127 -1119
rect -104 -1120 -78 -1116
rect -139 -1138 -127 -1134
rect -104 -1136 -101 -1120
rect -145 -1150 -141 -1146
rect -163 -1154 -141 -1150
rect -163 -1165 -156 -1154
rect -145 -1157 -141 -1154
rect -131 -1165 -127 -1138
rect -269 -1198 -253 -1194
rect -249 -1190 -231 -1186
rect -269 -1215 -265 -1198
rect -269 -1219 -258 -1215
rect -269 -1247 -264 -1219
rect -258 -1238 -252 -1227
rect -249 -1239 -246 -1190
rect -190 -1191 -187 -1169
rect -173 -1170 -156 -1165
rect -139 -1169 -127 -1165
rect -243 -1198 -195 -1194
rect -243 -1216 -240 -1198
rect -218 -1219 -206 -1215
rect -224 -1231 -220 -1227
rect -242 -1235 -220 -1231
rect -242 -1246 -235 -1235
rect -224 -1238 -220 -1235
rect -210 -1246 -206 -1219
rect -269 -1260 -262 -1247
rect -252 -1251 -235 -1246
rect -218 -1250 -206 -1246
rect -268 -1325 -262 -1260
rect -209 -1259 -206 -1250
rect -209 -1311 -205 -1259
rect -202 -1301 -195 -1198
rect -190 -1195 -179 -1191
rect -190 -1273 -185 -1195
rect -179 -1214 -173 -1203
rect -170 -1215 -167 -1170
rect -164 -1192 -161 -1170
rect -130 -1191 -127 -1169
rect -109 -1140 -101 -1136
rect -98 -1139 -90 -1135
rect -109 -1179 -106 -1140
rect -98 -1170 -95 -1139
rect -90 -1158 -84 -1147
rect -81 -1159 -78 -1120
rect -75 -1120 -20 -1116
rect 6 -1120 9 -1077
rect -75 -1136 -72 -1120
rect -50 -1139 -38 -1135
rect -56 -1151 -52 -1147
rect -74 -1155 -52 -1151
rect -74 -1166 -67 -1155
rect -56 -1158 -52 -1155
rect -42 -1166 -38 -1139
rect -84 -1171 -67 -1166
rect -50 -1170 -38 -1166
rect -109 -1182 -101 -1179
rect -73 -1182 -70 -1171
rect -41 -1179 -38 -1170
rect -29 -1182 -26 -1175
rect -139 -1195 -127 -1191
rect -145 -1207 -141 -1203
rect -163 -1211 -141 -1207
rect -163 -1222 -156 -1211
rect -145 -1214 -141 -1211
rect -131 -1222 -127 -1195
rect -173 -1227 -156 -1222
rect -139 -1226 -127 -1222
rect -162 -1251 -157 -1227
rect -124 -1202 -113 -1198
rect -124 -1232 -119 -1202
rect -113 -1221 -107 -1210
rect -104 -1222 -101 -1182
rect -98 -1187 -26 -1182
rect -98 -1199 -95 -1187
rect -49 -1194 -38 -1190
rect -73 -1202 -61 -1198
rect -79 -1214 -75 -1210
rect -97 -1218 -75 -1214
rect -97 -1229 -90 -1218
rect -79 -1221 -75 -1218
rect -65 -1229 -61 -1202
rect -49 -1225 -44 -1194
rect -38 -1213 -32 -1202
rect -29 -1214 -26 -1187
rect -23 -1191 -20 -1120
rect 7 -1126 9 -1120
rect 6 -1161 9 -1126
rect 76 -1082 144 -1072
rect 76 -1153 82 -1082
rect 161 -1094 168 -1063
rect 90 -1101 168 -1094
rect 214 -1090 220 -1058
rect 231 -1060 237 -1041
rect 264 -1049 267 -1040
rect 306 -1053 311 -1033
rect 339 -1042 342 -1032
rect 340 -1049 342 -1042
rect 275 -1059 311 -1053
rect 231 -1066 272 -1060
rect 249 -1075 260 -1071
rect 249 -1090 254 -1075
rect 214 -1096 254 -1090
rect 90 -1140 98 -1101
rect 249 -1106 254 -1096
rect 260 -1094 266 -1083
rect 269 -1095 272 -1066
rect 275 -1072 278 -1059
rect 300 -1075 312 -1071
rect 294 -1087 298 -1083
rect 276 -1091 298 -1087
rect 276 -1102 283 -1091
rect 294 -1094 298 -1091
rect 308 -1091 312 -1075
rect 339 -1091 342 -1049
rect 308 -1096 342 -1091
rect 308 -1102 312 -1096
rect 266 -1107 283 -1102
rect 300 -1106 312 -1102
rect 276 -1110 283 -1107
rect 163 -1117 283 -1110
rect 309 -1115 312 -1106
rect 137 -1129 147 -1120
rect 92 -1145 97 -1140
rect 142 -1141 147 -1129
rect 92 -1148 107 -1145
rect 76 -1156 88 -1153
rect 77 -1157 88 -1156
rect 6 -1165 14 -1161
rect 11 -1190 14 -1165
rect 2 -1194 14 -1190
rect -4 -1206 0 -1202
rect -22 -1210 0 -1206
rect -22 -1221 -15 -1210
rect -4 -1213 0 -1210
rect 10 -1221 14 -1194
rect 77 -1188 82 -1157
rect 88 -1176 94 -1165
rect 97 -1177 100 -1148
rect 103 -1150 107 -1148
rect 103 -1154 106 -1150
rect 143 -1153 146 -1141
rect 128 -1157 140 -1153
rect 122 -1169 126 -1165
rect 104 -1173 126 -1169
rect 104 -1184 111 -1173
rect 122 -1176 126 -1173
rect 136 -1184 140 -1157
rect 77 -1213 80 -1188
rect 94 -1189 111 -1184
rect 128 -1188 140 -1184
rect 98 -1205 102 -1189
rect 136 -1200 140 -1188
rect 139 -1205 140 -1200
rect 143 -1157 154 -1153
rect 143 -1188 148 -1157
rect 154 -1176 160 -1165
rect 163 -1177 166 -1117
rect 169 -1131 237 -1128
rect 169 -1154 172 -1131
rect 229 -1135 237 -1131
rect 276 -1135 283 -1117
rect 203 -1138 206 -1137
rect 201 -1153 206 -1138
rect 229 -1139 255 -1135
rect 194 -1157 206 -1153
rect 229 -1155 232 -1139
rect 188 -1169 192 -1165
rect 170 -1173 192 -1169
rect 170 -1184 177 -1173
rect 188 -1176 192 -1173
rect 202 -1184 206 -1157
rect -32 -1226 -15 -1221
rect 2 -1225 14 -1221
rect -124 -1238 -118 -1232
rect -107 -1234 -90 -1229
rect -73 -1233 -61 -1229
rect -124 -1242 -102 -1238
rect -162 -1254 -147 -1251
rect -177 -1263 -166 -1259
rect -177 -1273 -172 -1263
rect -190 -1277 -172 -1273
rect -177 -1294 -172 -1277
rect -166 -1282 -160 -1271
rect -157 -1283 -154 -1254
rect -151 -1256 -147 -1254
rect -151 -1260 -148 -1256
rect -126 -1263 -114 -1259
rect -132 -1275 -128 -1271
rect -150 -1279 -128 -1275
rect -150 -1290 -143 -1279
rect -132 -1282 -128 -1279
rect -118 -1290 -114 -1263
rect -160 -1295 -143 -1290
rect -126 -1294 -114 -1290
rect -154 -1301 -147 -1295
rect -202 -1307 -147 -1301
rect -154 -1308 -147 -1307
rect -117 -1311 -114 -1294
rect -209 -1316 -114 -1311
rect -108 -1325 -102 -1242
rect -97 -1253 -91 -1234
rect -64 -1242 -61 -1233
rect -22 -1246 -17 -1226
rect 11 -1234 14 -1225
rect 12 -1241 14 -1234
rect -53 -1252 -17 -1246
rect -97 -1256 -56 -1253
rect -92 -1259 -56 -1256
rect -79 -1268 -68 -1264
rect -79 -1299 -74 -1268
rect -68 -1287 -62 -1276
rect -59 -1288 -56 -1259
rect -53 -1265 -50 -1252
rect 11 -1264 14 -1241
rect -28 -1268 14 -1264
rect -20 -1269 14 -1268
rect 64 -1217 80 -1213
rect 84 -1209 102 -1205
rect 64 -1234 68 -1217
rect 64 -1238 75 -1234
rect 64 -1266 69 -1238
rect 75 -1257 81 -1246
rect 84 -1258 87 -1209
rect 143 -1210 146 -1188
rect 160 -1189 177 -1184
rect 194 -1188 206 -1184
rect 90 -1217 138 -1213
rect 90 -1235 93 -1217
rect 115 -1238 127 -1234
rect 109 -1250 113 -1246
rect 91 -1254 113 -1250
rect 91 -1265 98 -1254
rect 109 -1257 113 -1254
rect 123 -1265 127 -1238
rect -34 -1280 -30 -1276
rect -52 -1284 -30 -1280
rect -52 -1295 -45 -1284
rect -34 -1287 -30 -1284
rect -20 -1279 -17 -1269
rect 64 -1279 71 -1266
rect 81 -1270 98 -1265
rect 115 -1269 127 -1265
rect -20 -1295 -16 -1279
rect -79 -1325 -73 -1299
rect -62 -1300 -45 -1295
rect -28 -1299 -16 -1295
rect -268 -1333 -73 -1325
rect -268 -1334 -74 -1333
rect -229 -1348 -72 -1340
rect -79 -1352 -72 -1348
rect -80 -1378 -72 -1352
rect -59 -1402 -53 -1300
rect -19 -1308 -16 -1299
rect 65 -1344 71 -1279
rect 124 -1278 127 -1269
rect 124 -1330 128 -1278
rect 131 -1320 138 -1217
rect 143 -1214 154 -1210
rect 143 -1292 148 -1214
rect 154 -1233 160 -1222
rect 163 -1234 166 -1189
rect 169 -1211 172 -1189
rect 203 -1210 206 -1188
rect 224 -1159 232 -1155
rect 235 -1158 243 -1154
rect 224 -1198 227 -1159
rect 235 -1189 238 -1158
rect 243 -1177 249 -1166
rect 252 -1178 255 -1139
rect 258 -1139 313 -1135
rect 339 -1139 342 -1096
rect 681 -1009 684 -962
rect 681 -1013 692 -1009
rect 681 -1044 686 -1013
rect 692 -1032 698 -1021
rect 701 -1033 704 -954
rect 767 -963 784 -962
rect 799 -962 804 -954
rect 789 -963 793 -962
rect 767 -966 793 -963
rect 767 -982 770 -966
rect 707 -987 770 -982
rect 707 -1010 710 -987
rect 741 -1009 744 -993
rect 767 -1003 770 -987
rect 732 -1013 744 -1009
rect 726 -1025 730 -1021
rect 708 -1029 730 -1025
rect 708 -1040 715 -1029
rect 726 -1032 730 -1029
rect 740 -1040 744 -1013
rect 681 -1066 684 -1044
rect 698 -1045 715 -1040
rect 732 -1044 744 -1040
rect 753 -1044 757 -1003
rect 763 -1006 770 -1003
rect 773 -985 781 -981
rect 763 -1018 766 -1006
rect 773 -1009 776 -985
rect 781 -1004 787 -993
rect 790 -1005 793 -966
rect 796 -966 851 -962
rect 796 -982 799 -966
rect 821 -985 833 -981
rect 815 -997 819 -993
rect 797 -1001 819 -997
rect 797 -1012 804 -1001
rect 815 -1004 819 -1001
rect 829 -1012 833 -985
rect 787 -1017 804 -1012
rect 821 -1016 833 -1012
rect 763 -1022 770 -1018
rect 765 -1024 770 -1022
rect 681 -1070 692 -1066
rect 681 -1101 686 -1070
rect 692 -1089 698 -1078
rect 701 -1090 704 -1045
rect 707 -1067 710 -1045
rect 741 -1066 744 -1044
rect 732 -1070 744 -1066
rect 726 -1082 730 -1078
rect 708 -1086 730 -1082
rect 708 -1097 715 -1086
rect 726 -1089 730 -1086
rect 740 -1097 744 -1070
rect 748 -1048 758 -1044
rect 748 -1092 752 -1048
rect 758 -1067 764 -1056
rect 767 -1068 770 -1024
rect 798 -1028 801 -1017
rect 830 -1025 833 -1016
rect 773 -1033 845 -1028
rect 773 -1045 776 -1033
rect 822 -1040 833 -1036
rect 798 -1048 810 -1044
rect 792 -1060 796 -1056
rect 774 -1064 796 -1060
rect 774 -1075 781 -1064
rect 792 -1067 796 -1064
rect 806 -1075 810 -1048
rect 822 -1071 827 -1040
rect 833 -1059 839 -1048
rect 842 -1060 845 -1033
rect 848 -1037 851 -966
rect 880 -1036 885 -1011
rect 873 -1040 885 -1036
rect 867 -1052 871 -1048
rect 849 -1056 871 -1052
rect 849 -1067 856 -1056
rect 867 -1059 871 -1056
rect 881 -1067 885 -1040
rect 839 -1072 856 -1067
rect 873 -1071 885 -1067
rect 764 -1080 781 -1075
rect 798 -1079 810 -1075
rect 748 -1097 762 -1092
rect 682 -1111 686 -1101
rect 698 -1102 715 -1097
rect 732 -1101 744 -1097
rect 258 -1155 261 -1139
rect 283 -1158 295 -1154
rect 277 -1170 281 -1166
rect 259 -1174 281 -1170
rect 259 -1185 266 -1174
rect 277 -1177 281 -1174
rect 291 -1185 295 -1158
rect 249 -1190 266 -1185
rect 283 -1189 295 -1185
rect 224 -1201 232 -1198
rect 260 -1201 263 -1190
rect 292 -1198 295 -1189
rect 304 -1201 307 -1194
rect 194 -1214 206 -1210
rect 188 -1226 192 -1222
rect 170 -1230 192 -1226
rect 170 -1241 177 -1230
rect 188 -1233 192 -1230
rect 202 -1241 206 -1214
rect 160 -1246 177 -1241
rect 194 -1245 206 -1241
rect 171 -1270 176 -1246
rect 209 -1221 220 -1217
rect 209 -1251 214 -1221
rect 220 -1240 226 -1229
rect 229 -1241 232 -1201
rect 235 -1206 307 -1201
rect 235 -1218 238 -1206
rect 284 -1213 295 -1209
rect 260 -1221 272 -1217
rect 254 -1233 258 -1229
rect 236 -1237 258 -1233
rect 236 -1248 243 -1237
rect 254 -1240 258 -1237
rect 268 -1248 272 -1221
rect 284 -1244 289 -1213
rect 295 -1232 301 -1221
rect 304 -1233 307 -1206
rect 310 -1210 313 -1139
rect 340 -1145 342 -1139
rect 339 -1180 342 -1145
rect 619 -1121 687 -1111
rect 339 -1184 347 -1180
rect 344 -1209 347 -1184
rect 619 -1192 625 -1121
rect 704 -1133 711 -1102
rect 633 -1140 711 -1133
rect 757 -1129 763 -1097
rect 774 -1099 780 -1080
rect 807 -1088 810 -1079
rect 849 -1092 854 -1072
rect 882 -1081 885 -1071
rect 883 -1088 885 -1081
rect 818 -1098 854 -1092
rect 774 -1105 815 -1099
rect 792 -1114 803 -1110
rect 792 -1129 797 -1114
rect 757 -1135 797 -1129
rect 633 -1179 641 -1140
rect 792 -1145 797 -1135
rect 803 -1133 809 -1122
rect 812 -1134 815 -1105
rect 818 -1111 821 -1098
rect 843 -1114 855 -1110
rect 837 -1126 841 -1122
rect 819 -1130 841 -1126
rect 819 -1141 826 -1130
rect 837 -1133 841 -1130
rect 851 -1130 855 -1114
rect 882 -1130 885 -1088
rect 851 -1135 885 -1130
rect 851 -1141 855 -1135
rect 809 -1146 826 -1141
rect 843 -1145 855 -1141
rect 819 -1149 826 -1146
rect 706 -1156 826 -1149
rect 852 -1154 855 -1145
rect 680 -1168 690 -1159
rect 635 -1184 640 -1179
rect 685 -1180 690 -1168
rect 635 -1187 650 -1184
rect 619 -1195 631 -1192
rect 335 -1213 347 -1209
rect 329 -1225 333 -1221
rect 311 -1229 333 -1225
rect 311 -1240 318 -1229
rect 329 -1232 333 -1229
rect 343 -1240 347 -1213
rect 301 -1245 318 -1240
rect 335 -1244 347 -1240
rect 209 -1257 215 -1251
rect 226 -1253 243 -1248
rect 260 -1252 272 -1248
rect 209 -1261 231 -1257
rect 171 -1273 186 -1270
rect 156 -1282 167 -1278
rect 156 -1292 161 -1282
rect 143 -1296 161 -1292
rect 156 -1313 161 -1296
rect 167 -1301 173 -1290
rect 176 -1302 179 -1273
rect 182 -1275 186 -1273
rect 182 -1279 185 -1275
rect 207 -1282 219 -1278
rect 201 -1294 205 -1290
rect 183 -1298 205 -1294
rect 183 -1309 190 -1298
rect 201 -1301 205 -1298
rect 215 -1309 219 -1282
rect 173 -1314 190 -1309
rect 207 -1313 219 -1309
rect 179 -1320 186 -1314
rect 131 -1326 186 -1320
rect 179 -1327 186 -1326
rect 216 -1330 219 -1313
rect 124 -1335 219 -1330
rect 225 -1344 231 -1261
rect 236 -1272 242 -1253
rect 269 -1261 272 -1252
rect 311 -1265 316 -1245
rect 344 -1253 347 -1244
rect 620 -1196 631 -1195
rect 620 -1227 625 -1196
rect 631 -1215 637 -1204
rect 640 -1216 643 -1187
rect 646 -1189 650 -1187
rect 646 -1193 649 -1189
rect 686 -1192 689 -1180
rect 671 -1196 683 -1192
rect 665 -1208 669 -1204
rect 647 -1212 669 -1208
rect 647 -1223 654 -1212
rect 665 -1215 669 -1212
rect 679 -1223 683 -1196
rect 620 -1252 623 -1227
rect 637 -1228 654 -1223
rect 671 -1227 683 -1223
rect 641 -1244 645 -1228
rect 679 -1239 683 -1227
rect 682 -1244 683 -1239
rect 686 -1196 697 -1192
rect 686 -1227 691 -1196
rect 697 -1215 703 -1204
rect 706 -1216 709 -1156
rect 712 -1170 780 -1167
rect 712 -1193 715 -1170
rect 772 -1174 780 -1170
rect 819 -1174 826 -1156
rect 746 -1177 749 -1176
rect 744 -1192 749 -1177
rect 772 -1178 798 -1174
rect 737 -1196 749 -1192
rect 772 -1194 775 -1178
rect 731 -1208 735 -1204
rect 713 -1212 735 -1208
rect 713 -1223 720 -1212
rect 731 -1215 735 -1212
rect 745 -1223 749 -1196
rect 345 -1260 347 -1253
rect 280 -1271 316 -1265
rect 236 -1275 277 -1272
rect 241 -1278 277 -1275
rect 254 -1287 265 -1283
rect 254 -1318 259 -1287
rect 265 -1306 271 -1295
rect 274 -1307 277 -1278
rect 280 -1284 283 -1271
rect 344 -1283 347 -1260
rect 305 -1287 347 -1283
rect 313 -1288 347 -1287
rect 607 -1256 623 -1252
rect 627 -1248 645 -1244
rect 607 -1273 611 -1256
rect 607 -1277 618 -1273
rect 299 -1299 303 -1295
rect 281 -1303 303 -1299
rect 281 -1314 288 -1303
rect 299 -1306 303 -1303
rect 313 -1314 317 -1288
rect 254 -1344 260 -1318
rect 271 -1319 288 -1314
rect 305 -1318 317 -1314
rect 607 -1305 612 -1277
rect 618 -1296 624 -1285
rect 627 -1297 630 -1248
rect 686 -1249 689 -1227
rect 703 -1228 720 -1223
rect 737 -1227 749 -1223
rect 633 -1256 681 -1252
rect 633 -1274 636 -1256
rect 658 -1277 670 -1273
rect 652 -1289 656 -1285
rect 634 -1293 656 -1289
rect 634 -1304 641 -1293
rect 652 -1296 656 -1293
rect 666 -1304 670 -1277
rect 607 -1318 614 -1305
rect 624 -1309 641 -1304
rect 658 -1308 670 -1304
rect 65 -1352 260 -1344
rect 65 -1353 259 -1352
rect 69 -1380 76 -1353
rect 104 -1367 261 -1359
rect 189 -1380 197 -1376
rect 70 -1387 197 -1380
rect -59 -1408 182 -1402
rect -373 -1456 -363 -1426
rect -281 -1432 153 -1425
rect -373 -1463 -185 -1456
rect -162 -1463 -14 -1456
rect -463 -1509 -380 -1500
rect -462 -1542 -457 -1509
rect -388 -1510 -380 -1509
rect -350 -1538 -347 -1537
rect -462 -1546 -456 -1542
rect -498 -1558 -492 -1547
rect -461 -1556 -456 -1546
rect -449 -1543 -347 -1538
rect -449 -1577 -443 -1543
rect -544 -1581 -440 -1577
rect -564 -1636 -561 -1589
rect -564 -1640 -553 -1636
rect -564 -1671 -559 -1640
rect -553 -1659 -547 -1648
rect -544 -1660 -541 -1581
rect -478 -1590 -461 -1589
rect -446 -1589 -441 -1581
rect -456 -1590 -452 -1589
rect -478 -1593 -452 -1590
rect -478 -1609 -475 -1593
rect -538 -1614 -475 -1609
rect -538 -1637 -535 -1614
rect -504 -1636 -501 -1620
rect -478 -1630 -475 -1614
rect -513 -1640 -501 -1636
rect -519 -1652 -515 -1648
rect -537 -1656 -515 -1652
rect -537 -1667 -530 -1656
rect -519 -1659 -515 -1656
rect -505 -1667 -501 -1640
rect -564 -1693 -561 -1671
rect -547 -1672 -530 -1667
rect -513 -1671 -501 -1667
rect -492 -1671 -488 -1630
rect -482 -1633 -475 -1630
rect -472 -1612 -464 -1608
rect -482 -1645 -479 -1633
rect -472 -1636 -469 -1612
rect -464 -1631 -458 -1620
rect -455 -1632 -452 -1593
rect -449 -1593 -394 -1589
rect -449 -1609 -446 -1593
rect -424 -1612 -412 -1608
rect -430 -1624 -426 -1620
rect -448 -1628 -426 -1624
rect -448 -1639 -441 -1628
rect -430 -1631 -426 -1628
rect -416 -1639 -412 -1612
rect -458 -1644 -441 -1639
rect -424 -1643 -412 -1639
rect -482 -1649 -475 -1645
rect -480 -1651 -475 -1649
rect -564 -1697 -553 -1693
rect -564 -1728 -559 -1697
rect -553 -1716 -547 -1705
rect -544 -1717 -541 -1672
rect -538 -1694 -535 -1672
rect -504 -1693 -501 -1671
rect -513 -1697 -501 -1693
rect -519 -1709 -515 -1705
rect -537 -1713 -515 -1709
rect -537 -1724 -530 -1713
rect -519 -1716 -515 -1713
rect -505 -1724 -501 -1697
rect -497 -1675 -487 -1671
rect -497 -1719 -493 -1675
rect -487 -1694 -481 -1683
rect -478 -1695 -475 -1651
rect -447 -1655 -444 -1644
rect -415 -1652 -412 -1643
rect -472 -1660 -400 -1655
rect -472 -1672 -469 -1660
rect -423 -1667 -412 -1663
rect -447 -1675 -435 -1671
rect -453 -1687 -449 -1683
rect -471 -1691 -449 -1687
rect -471 -1702 -464 -1691
rect -453 -1694 -449 -1691
rect -439 -1702 -435 -1675
rect -423 -1698 -418 -1667
rect -412 -1686 -406 -1675
rect -403 -1687 -400 -1660
rect -397 -1664 -394 -1593
rect -365 -1663 -360 -1638
rect -372 -1667 -360 -1663
rect -378 -1679 -374 -1675
rect -396 -1683 -374 -1679
rect -396 -1694 -389 -1683
rect -378 -1686 -374 -1683
rect -364 -1694 -360 -1667
rect -406 -1699 -389 -1694
rect -372 -1698 -360 -1694
rect -481 -1707 -464 -1702
rect -447 -1706 -435 -1702
rect -497 -1724 -483 -1719
rect -563 -1738 -559 -1728
rect -547 -1729 -530 -1724
rect -513 -1728 -501 -1724
rect -626 -1748 -558 -1738
rect -626 -1819 -620 -1748
rect -541 -1760 -534 -1729
rect -612 -1767 -534 -1760
rect -488 -1756 -482 -1724
rect -471 -1726 -465 -1707
rect -438 -1715 -435 -1706
rect -396 -1719 -391 -1699
rect -363 -1708 -360 -1698
rect -362 -1715 -360 -1708
rect -427 -1725 -391 -1719
rect -471 -1732 -430 -1726
rect -453 -1741 -442 -1737
rect -453 -1756 -448 -1741
rect -488 -1762 -448 -1756
rect -612 -1806 -604 -1767
rect -453 -1772 -448 -1762
rect -442 -1760 -436 -1749
rect -433 -1761 -430 -1732
rect -427 -1738 -424 -1725
rect -402 -1741 -390 -1737
rect -408 -1753 -404 -1749
rect -426 -1757 -404 -1753
rect -426 -1768 -419 -1757
rect -408 -1760 -404 -1757
rect -394 -1757 -390 -1741
rect -363 -1757 -360 -1715
rect -394 -1762 -360 -1757
rect -394 -1768 -390 -1762
rect -436 -1773 -419 -1768
rect -402 -1772 -390 -1768
rect -426 -1776 -419 -1773
rect -539 -1783 -419 -1776
rect -393 -1781 -390 -1772
rect -565 -1795 -555 -1786
rect -610 -1811 -605 -1806
rect -560 -1807 -555 -1795
rect -610 -1814 -595 -1811
rect -626 -1822 -614 -1819
rect -625 -1823 -614 -1822
rect -625 -1854 -620 -1823
rect -614 -1842 -608 -1831
rect -605 -1843 -602 -1814
rect -599 -1816 -595 -1814
rect -599 -1820 -596 -1816
rect -559 -1819 -556 -1807
rect -574 -1823 -562 -1819
rect -580 -1835 -576 -1831
rect -598 -1839 -576 -1835
rect -598 -1850 -591 -1839
rect -580 -1842 -576 -1839
rect -566 -1850 -562 -1823
rect -625 -1879 -622 -1854
rect -608 -1855 -591 -1850
rect -574 -1854 -562 -1850
rect -604 -1871 -600 -1855
rect -566 -1866 -562 -1854
rect -563 -1871 -562 -1866
rect -559 -1823 -548 -1819
rect -559 -1854 -554 -1823
rect -548 -1842 -542 -1831
rect -539 -1843 -536 -1783
rect -533 -1797 -465 -1794
rect -533 -1820 -530 -1797
rect -473 -1801 -465 -1797
rect -426 -1801 -419 -1783
rect -499 -1804 -496 -1803
rect -501 -1819 -496 -1804
rect -473 -1805 -447 -1801
rect -508 -1823 -496 -1819
rect -473 -1821 -470 -1805
rect -514 -1835 -510 -1831
rect -532 -1839 -510 -1835
rect -532 -1850 -525 -1839
rect -514 -1842 -510 -1839
rect -500 -1850 -496 -1823
rect -638 -1883 -622 -1879
rect -618 -1875 -600 -1871
rect -638 -1900 -634 -1883
rect -638 -1904 -627 -1900
rect -638 -1932 -633 -1904
rect -627 -1923 -621 -1912
rect -618 -1924 -615 -1875
rect -559 -1876 -556 -1854
rect -542 -1855 -525 -1850
rect -508 -1854 -496 -1850
rect -612 -1883 -564 -1879
rect -612 -1901 -609 -1883
rect -587 -1904 -575 -1900
rect -593 -1916 -589 -1912
rect -611 -1920 -589 -1916
rect -611 -1931 -604 -1920
rect -593 -1923 -589 -1920
rect -579 -1931 -575 -1904
rect -638 -1945 -631 -1932
rect -621 -1936 -604 -1931
rect -587 -1935 -575 -1931
rect -637 -2010 -631 -1945
rect -578 -1944 -575 -1935
rect -578 -1996 -574 -1944
rect -571 -1986 -564 -1883
rect -559 -1880 -548 -1876
rect -559 -1958 -554 -1880
rect -548 -1899 -542 -1888
rect -539 -1900 -536 -1855
rect -533 -1877 -530 -1855
rect -499 -1876 -496 -1854
rect -478 -1825 -470 -1821
rect -467 -1824 -459 -1820
rect -478 -1864 -475 -1825
rect -467 -1855 -464 -1824
rect -459 -1843 -453 -1832
rect -450 -1844 -447 -1805
rect -444 -1805 -389 -1801
rect -363 -1805 -360 -1762
rect -444 -1821 -441 -1805
rect -419 -1824 -407 -1820
rect -425 -1836 -421 -1832
rect -443 -1840 -421 -1836
rect -443 -1851 -436 -1840
rect -425 -1843 -421 -1840
rect -411 -1851 -407 -1824
rect -453 -1856 -436 -1851
rect -419 -1855 -407 -1851
rect -478 -1867 -470 -1864
rect -442 -1867 -439 -1856
rect -410 -1864 -407 -1855
rect -398 -1867 -395 -1860
rect -508 -1880 -496 -1876
rect -514 -1892 -510 -1888
rect -532 -1896 -510 -1892
rect -532 -1907 -525 -1896
rect -514 -1899 -510 -1896
rect -500 -1907 -496 -1880
rect -542 -1912 -525 -1907
rect -508 -1911 -496 -1907
rect -531 -1936 -526 -1912
rect -493 -1887 -482 -1883
rect -493 -1917 -488 -1887
rect -482 -1906 -476 -1895
rect -473 -1907 -470 -1867
rect -467 -1872 -395 -1867
rect -467 -1884 -464 -1872
rect -418 -1879 -407 -1875
rect -442 -1887 -430 -1883
rect -448 -1899 -444 -1895
rect -466 -1903 -444 -1899
rect -466 -1914 -459 -1903
rect -448 -1906 -444 -1903
rect -434 -1914 -430 -1887
rect -418 -1910 -413 -1879
rect -407 -1898 -401 -1887
rect -398 -1899 -395 -1872
rect -392 -1876 -389 -1805
rect -362 -1811 -360 -1805
rect -363 -1846 -360 -1811
rect -363 -1850 -355 -1846
rect -358 -1875 -355 -1850
rect -367 -1879 -355 -1875
rect -373 -1891 -369 -1887
rect -391 -1895 -369 -1891
rect -391 -1906 -384 -1895
rect -373 -1898 -369 -1895
rect -359 -1906 -355 -1879
rect -401 -1911 -384 -1906
rect -367 -1910 -355 -1906
rect -493 -1923 -487 -1917
rect -476 -1919 -459 -1914
rect -442 -1918 -430 -1914
rect -493 -1927 -471 -1923
rect -531 -1939 -516 -1936
rect -546 -1948 -535 -1944
rect -546 -1958 -541 -1948
rect -559 -1962 -541 -1958
rect -546 -1979 -541 -1962
rect -535 -1967 -529 -1956
rect -526 -1968 -523 -1939
rect -520 -1941 -516 -1939
rect -520 -1945 -517 -1941
rect -495 -1948 -483 -1944
rect -501 -1960 -497 -1956
rect -519 -1964 -497 -1960
rect -519 -1975 -512 -1964
rect -501 -1967 -497 -1964
rect -487 -1975 -483 -1948
rect -529 -1980 -512 -1975
rect -495 -1979 -483 -1975
rect -523 -1986 -516 -1980
rect -571 -1992 -516 -1986
rect -523 -1993 -516 -1992
rect -486 -1996 -483 -1979
rect -578 -2001 -483 -1996
rect -477 -2010 -471 -1927
rect -466 -1938 -460 -1919
rect -433 -1927 -430 -1918
rect -391 -1931 -386 -1911
rect -358 -1919 -355 -1910
rect -357 -1926 -355 -1919
rect -422 -1937 -386 -1931
rect -466 -1941 -425 -1938
rect -461 -1944 -425 -1941
rect -448 -1953 -437 -1949
rect -448 -1984 -443 -1953
rect -437 -1972 -431 -1961
rect -428 -1973 -425 -1944
rect -422 -1950 -419 -1937
rect -358 -1949 -355 -1926
rect -397 -1953 -355 -1949
rect -389 -1954 -355 -1953
rect -403 -1965 -399 -1961
rect -421 -1969 -399 -1965
rect -421 -1980 -414 -1969
rect -403 -1972 -399 -1969
rect -389 -1980 -385 -1954
rect -448 -2010 -442 -1984
rect -431 -1985 -414 -1980
rect -397 -1984 -385 -1980
rect -637 -2018 -442 -2010
rect -637 -2019 -443 -2018
rect -598 -2033 -441 -2025
rect -448 -2252 -441 -2033
rect -449 -2263 -441 -2252
rect -428 -2263 -422 -1985
rect -388 -1993 -385 -1984
rect -350 -1994 -347 -1543
rect -259 -1580 -256 -1476
rect -193 -1477 -185 -1463
rect -193 -1488 -186 -1477
rect -157 -1487 -151 -1463
rect -193 -1502 -187 -1488
rect -156 -1500 -151 -1487
rect -145 -1476 -31 -1470
rect -145 -1484 -138 -1476
rect -145 -1487 -137 -1484
rect -145 -1521 -138 -1487
rect -239 -1525 -135 -1521
rect -259 -1584 -248 -1580
rect -259 -1615 -254 -1584
rect -248 -1603 -242 -1592
rect -239 -1604 -236 -1525
rect -173 -1534 -156 -1533
rect -141 -1533 -136 -1525
rect -151 -1534 -147 -1533
rect -173 -1537 -147 -1534
rect -173 -1553 -170 -1537
rect -233 -1558 -170 -1553
rect -233 -1581 -230 -1558
rect -199 -1580 -196 -1564
rect -173 -1574 -170 -1558
rect -208 -1584 -196 -1580
rect -214 -1596 -210 -1592
rect -232 -1600 -210 -1596
rect -232 -1611 -225 -1600
rect -214 -1603 -210 -1600
rect -200 -1611 -196 -1584
rect -259 -1637 -256 -1615
rect -242 -1616 -225 -1611
rect -208 -1615 -196 -1611
rect -187 -1615 -183 -1574
rect -177 -1577 -170 -1574
rect -167 -1556 -159 -1552
rect -177 -1589 -174 -1577
rect -167 -1580 -164 -1556
rect -159 -1575 -153 -1564
rect -150 -1576 -147 -1537
rect -144 -1537 -89 -1533
rect -144 -1553 -141 -1537
rect -119 -1556 -107 -1552
rect -125 -1568 -121 -1564
rect -143 -1572 -121 -1568
rect -143 -1583 -136 -1572
rect -125 -1575 -121 -1572
rect -111 -1583 -107 -1556
rect -153 -1588 -136 -1583
rect -119 -1587 -107 -1583
rect -177 -1593 -170 -1589
rect -175 -1595 -170 -1593
rect -259 -1641 -248 -1637
rect -259 -1672 -254 -1641
rect -248 -1660 -242 -1649
rect -239 -1661 -236 -1616
rect -233 -1638 -230 -1616
rect -199 -1637 -196 -1615
rect -208 -1641 -196 -1637
rect -214 -1653 -210 -1649
rect -232 -1657 -210 -1653
rect -232 -1668 -225 -1657
rect -214 -1660 -210 -1657
rect -200 -1668 -196 -1641
rect -192 -1619 -182 -1615
rect -192 -1663 -188 -1619
rect -182 -1638 -176 -1627
rect -173 -1639 -170 -1595
rect -142 -1599 -139 -1588
rect -110 -1596 -107 -1587
rect -167 -1604 -95 -1599
rect -167 -1616 -164 -1604
rect -118 -1611 -107 -1607
rect -142 -1619 -130 -1615
rect -148 -1631 -144 -1627
rect -166 -1635 -144 -1631
rect -166 -1646 -159 -1635
rect -148 -1638 -144 -1635
rect -134 -1646 -130 -1619
rect -118 -1642 -113 -1611
rect -107 -1630 -101 -1619
rect -98 -1631 -95 -1604
rect -92 -1608 -89 -1537
rect -60 -1607 -55 -1582
rect -67 -1611 -55 -1607
rect -73 -1623 -69 -1619
rect -91 -1627 -69 -1623
rect -91 -1638 -84 -1627
rect -73 -1630 -69 -1627
rect -59 -1638 -55 -1611
rect -101 -1643 -84 -1638
rect -67 -1642 -55 -1638
rect -176 -1651 -159 -1646
rect -142 -1650 -130 -1646
rect -192 -1668 -178 -1663
rect -258 -1682 -254 -1672
rect -242 -1673 -225 -1668
rect -208 -1672 -196 -1668
rect -321 -1692 -253 -1682
rect -321 -1763 -315 -1692
rect -236 -1704 -229 -1673
rect -307 -1711 -229 -1704
rect -183 -1700 -177 -1668
rect -166 -1670 -160 -1651
rect -133 -1659 -130 -1650
rect -91 -1663 -86 -1643
rect -58 -1652 -55 -1642
rect -57 -1659 -55 -1652
rect -122 -1669 -86 -1663
rect -166 -1676 -125 -1670
rect -148 -1685 -137 -1681
rect -148 -1700 -143 -1685
rect -183 -1706 -143 -1700
rect -307 -1750 -299 -1711
rect -148 -1716 -143 -1706
rect -137 -1704 -131 -1693
rect -128 -1705 -125 -1676
rect -122 -1682 -119 -1669
rect -97 -1685 -85 -1681
rect -103 -1697 -99 -1693
rect -121 -1701 -99 -1697
rect -121 -1712 -114 -1701
rect -103 -1704 -99 -1701
rect -89 -1701 -85 -1685
rect -58 -1701 -55 -1659
rect -89 -1706 -55 -1701
rect -89 -1712 -85 -1706
rect -131 -1717 -114 -1712
rect -97 -1716 -85 -1712
rect -121 -1720 -114 -1717
rect -234 -1727 -114 -1720
rect -88 -1725 -85 -1716
rect -260 -1739 -250 -1730
rect -305 -1755 -300 -1750
rect -255 -1751 -250 -1739
rect -305 -1758 -290 -1755
rect -321 -1766 -309 -1763
rect -320 -1767 -309 -1766
rect -320 -1798 -315 -1767
rect -309 -1786 -303 -1775
rect -300 -1787 -297 -1758
rect -294 -1760 -290 -1758
rect -294 -1764 -291 -1760
rect -254 -1763 -251 -1751
rect -269 -1767 -257 -1763
rect -275 -1779 -271 -1775
rect -293 -1783 -271 -1779
rect -293 -1794 -286 -1783
rect -275 -1786 -271 -1783
rect -261 -1794 -257 -1767
rect -320 -1823 -317 -1798
rect -303 -1799 -286 -1794
rect -269 -1798 -257 -1794
rect -299 -1815 -295 -1799
rect -261 -1810 -257 -1798
rect -258 -1815 -257 -1810
rect -254 -1767 -243 -1763
rect -254 -1798 -249 -1767
rect -243 -1786 -237 -1775
rect -234 -1787 -231 -1727
rect -228 -1741 -160 -1738
rect -228 -1764 -225 -1741
rect -168 -1745 -160 -1741
rect -121 -1745 -114 -1727
rect -194 -1748 -191 -1747
rect -196 -1763 -191 -1748
rect -168 -1749 -142 -1745
rect -203 -1767 -191 -1763
rect -168 -1765 -165 -1749
rect -209 -1779 -205 -1775
rect -227 -1783 -205 -1779
rect -227 -1794 -220 -1783
rect -209 -1786 -205 -1783
rect -195 -1794 -191 -1767
rect -333 -1827 -317 -1823
rect -313 -1819 -295 -1815
rect -333 -1844 -329 -1827
rect -333 -1848 -322 -1844
rect -333 -1876 -328 -1848
rect -322 -1867 -316 -1856
rect -313 -1868 -310 -1819
rect -254 -1820 -251 -1798
rect -237 -1799 -220 -1794
rect -203 -1798 -191 -1794
rect -307 -1827 -259 -1823
rect -307 -1845 -304 -1827
rect -282 -1848 -270 -1844
rect -288 -1860 -284 -1856
rect -306 -1864 -284 -1860
rect -306 -1875 -299 -1864
rect -288 -1867 -284 -1864
rect -274 -1875 -270 -1848
rect -333 -1889 -326 -1876
rect -316 -1880 -299 -1875
rect -282 -1879 -270 -1875
rect -332 -1954 -326 -1889
rect -273 -1888 -270 -1879
rect -273 -1940 -269 -1888
rect -266 -1930 -259 -1827
rect -254 -1824 -243 -1820
rect -254 -1902 -249 -1824
rect -243 -1843 -237 -1832
rect -234 -1844 -231 -1799
rect -228 -1821 -225 -1799
rect -194 -1820 -191 -1798
rect -173 -1769 -165 -1765
rect -162 -1768 -154 -1764
rect -173 -1808 -170 -1769
rect -162 -1799 -159 -1768
rect -154 -1787 -148 -1776
rect -145 -1788 -142 -1749
rect -139 -1749 -84 -1745
rect -58 -1749 -55 -1706
rect -139 -1765 -136 -1749
rect -114 -1768 -102 -1764
rect -120 -1780 -116 -1776
rect -138 -1784 -116 -1780
rect -138 -1795 -131 -1784
rect -120 -1787 -116 -1784
rect -106 -1795 -102 -1768
rect -148 -1800 -131 -1795
rect -114 -1799 -102 -1795
rect -173 -1811 -165 -1808
rect -137 -1811 -134 -1800
rect -105 -1808 -102 -1799
rect -93 -1811 -90 -1804
rect -203 -1824 -191 -1820
rect -209 -1836 -205 -1832
rect -227 -1840 -205 -1836
rect -227 -1851 -220 -1840
rect -209 -1843 -205 -1840
rect -195 -1851 -191 -1824
rect -237 -1856 -220 -1851
rect -203 -1855 -191 -1851
rect -226 -1880 -221 -1856
rect -188 -1831 -177 -1827
rect -188 -1861 -183 -1831
rect -177 -1850 -171 -1839
rect -168 -1851 -165 -1811
rect -162 -1816 -90 -1811
rect -162 -1828 -159 -1816
rect -113 -1823 -102 -1819
rect -137 -1831 -125 -1827
rect -143 -1843 -139 -1839
rect -161 -1847 -139 -1843
rect -161 -1858 -154 -1847
rect -143 -1850 -139 -1847
rect -129 -1858 -125 -1831
rect -113 -1854 -108 -1823
rect -102 -1842 -96 -1831
rect -93 -1843 -90 -1816
rect -87 -1820 -84 -1749
rect -57 -1755 -55 -1749
rect -58 -1790 -55 -1755
rect -58 -1794 -50 -1790
rect -53 -1819 -50 -1794
rect -62 -1823 -50 -1819
rect -68 -1835 -64 -1831
rect -86 -1839 -64 -1835
rect -86 -1850 -79 -1839
rect -68 -1842 -64 -1839
rect -54 -1850 -50 -1823
rect -96 -1855 -79 -1850
rect -62 -1854 -50 -1850
rect -188 -1867 -182 -1861
rect -171 -1863 -154 -1858
rect -137 -1862 -125 -1858
rect -188 -1871 -166 -1867
rect -226 -1883 -211 -1880
rect -241 -1892 -230 -1888
rect -241 -1902 -236 -1892
rect -254 -1906 -236 -1902
rect -241 -1923 -236 -1906
rect -230 -1911 -224 -1900
rect -221 -1912 -218 -1883
rect -215 -1885 -211 -1883
rect -215 -1889 -212 -1885
rect -190 -1892 -178 -1888
rect -196 -1904 -192 -1900
rect -214 -1908 -192 -1904
rect -214 -1919 -207 -1908
rect -196 -1911 -192 -1908
rect -182 -1919 -178 -1892
rect -224 -1924 -207 -1919
rect -190 -1923 -178 -1919
rect -218 -1930 -211 -1924
rect -266 -1936 -211 -1930
rect -218 -1937 -211 -1936
rect -181 -1940 -178 -1923
rect -273 -1945 -178 -1940
rect -172 -1954 -166 -1871
rect -161 -1882 -155 -1863
rect -128 -1871 -125 -1862
rect -86 -1875 -81 -1855
rect -53 -1863 -50 -1854
rect -52 -1870 -50 -1863
rect -117 -1881 -81 -1875
rect -161 -1885 -120 -1882
rect -156 -1888 -120 -1885
rect -143 -1897 -132 -1893
rect -143 -1928 -138 -1897
rect -132 -1916 -126 -1905
rect -123 -1917 -120 -1888
rect -117 -1894 -114 -1881
rect -53 -1893 -50 -1870
rect -92 -1897 -50 -1893
rect -84 -1898 -50 -1897
rect -98 -1909 -94 -1905
rect -116 -1913 -94 -1909
rect -116 -1924 -109 -1913
rect -98 -1916 -94 -1913
rect -84 -1924 -80 -1898
rect -143 -1954 -137 -1928
rect -126 -1929 -109 -1924
rect -92 -1928 -80 -1924
rect -332 -1962 -137 -1954
rect -332 -1963 -138 -1962
rect -293 -1977 -141 -1969
rect -148 -1981 -141 -1977
rect -149 -1994 -141 -1981
rect -350 -2001 -141 -1994
rect -149 -2014 -141 -2001
rect -123 -2277 -117 -1929
rect -83 -1937 -80 -1928
rect -35 -2030 -31 -1476
rect -22 -2014 -16 -1463
rect 146 -1499 153 -1432
rect 176 -1492 182 -1408
rect 189 -1449 197 -1387
rect 254 -1393 261 -1367
rect 274 -1428 280 -1319
rect 314 -1327 317 -1318
rect 608 -1383 614 -1318
rect 667 -1317 670 -1308
rect 667 -1369 671 -1317
rect 674 -1359 681 -1256
rect 686 -1253 697 -1249
rect 686 -1331 691 -1253
rect 697 -1272 703 -1261
rect 706 -1273 709 -1228
rect 712 -1250 715 -1228
rect 746 -1249 749 -1227
rect 767 -1198 775 -1194
rect 778 -1197 786 -1193
rect 767 -1237 770 -1198
rect 778 -1228 781 -1197
rect 786 -1216 792 -1205
rect 795 -1217 798 -1178
rect 801 -1178 856 -1174
rect 882 -1178 885 -1135
rect 801 -1194 804 -1178
rect 826 -1197 838 -1193
rect 820 -1209 824 -1205
rect 802 -1213 824 -1209
rect 802 -1224 809 -1213
rect 820 -1216 824 -1213
rect 834 -1224 838 -1197
rect 792 -1229 809 -1224
rect 826 -1228 838 -1224
rect 767 -1240 775 -1237
rect 803 -1240 806 -1229
rect 835 -1237 838 -1228
rect 847 -1240 850 -1233
rect 737 -1253 749 -1249
rect 731 -1265 735 -1261
rect 713 -1269 735 -1265
rect 713 -1280 720 -1269
rect 731 -1272 735 -1269
rect 745 -1280 749 -1253
rect 703 -1285 720 -1280
rect 737 -1284 749 -1280
rect 714 -1309 719 -1285
rect 752 -1260 763 -1256
rect 752 -1290 757 -1260
rect 763 -1279 769 -1268
rect 772 -1280 775 -1240
rect 778 -1245 850 -1240
rect 778 -1257 781 -1245
rect 827 -1252 838 -1248
rect 803 -1260 815 -1256
rect 797 -1272 801 -1268
rect 779 -1276 801 -1272
rect 779 -1287 786 -1276
rect 797 -1279 801 -1276
rect 811 -1287 815 -1260
rect 827 -1283 832 -1252
rect 838 -1271 844 -1260
rect 847 -1272 850 -1245
rect 853 -1249 856 -1178
rect 883 -1184 885 -1178
rect 882 -1219 885 -1184
rect 882 -1223 890 -1219
rect 887 -1248 890 -1223
rect 878 -1252 890 -1248
rect 872 -1264 876 -1260
rect 854 -1268 876 -1264
rect 854 -1279 861 -1268
rect 872 -1271 876 -1268
rect 886 -1279 890 -1252
rect 844 -1284 861 -1279
rect 878 -1283 890 -1279
rect 752 -1296 758 -1290
rect 769 -1292 786 -1287
rect 803 -1291 815 -1287
rect 752 -1300 774 -1296
rect 714 -1312 729 -1309
rect 699 -1321 710 -1317
rect 699 -1331 704 -1321
rect 686 -1335 704 -1331
rect 699 -1352 704 -1335
rect 710 -1340 716 -1329
rect 719 -1341 722 -1312
rect 725 -1314 729 -1312
rect 725 -1318 728 -1314
rect 750 -1321 762 -1317
rect 744 -1333 748 -1329
rect 726 -1337 748 -1333
rect 726 -1348 733 -1337
rect 744 -1340 748 -1337
rect 758 -1348 762 -1321
rect 716 -1353 733 -1348
rect 750 -1352 762 -1348
rect 722 -1359 729 -1353
rect 674 -1365 729 -1359
rect 722 -1366 729 -1365
rect 759 -1369 762 -1352
rect 667 -1374 762 -1369
rect 768 -1383 774 -1300
rect 779 -1311 785 -1292
rect 812 -1300 815 -1291
rect 854 -1304 859 -1284
rect 887 -1292 890 -1283
rect 888 -1299 890 -1292
rect 823 -1310 859 -1304
rect 779 -1314 820 -1311
rect 784 -1317 820 -1314
rect 797 -1326 808 -1322
rect 797 -1357 802 -1326
rect 808 -1345 814 -1334
rect 817 -1346 820 -1317
rect 823 -1323 826 -1310
rect 887 -1322 890 -1299
rect 848 -1326 890 -1322
rect 856 -1327 890 -1326
rect 842 -1338 846 -1334
rect 824 -1342 846 -1338
rect 824 -1353 831 -1342
rect 842 -1345 846 -1342
rect 856 -1353 860 -1327
rect 797 -1383 803 -1357
rect 814 -1358 831 -1353
rect 848 -1357 860 -1353
rect 608 -1391 803 -1383
rect 608 -1392 802 -1391
rect 647 -1406 804 -1398
rect 797 -1410 804 -1406
rect 274 -1434 493 -1428
rect 274 -1435 280 -1434
rect 384 -1449 388 -1447
rect 189 -1454 388 -1449
rect 486 -1444 493 -1434
rect 796 -1437 804 -1410
rect 487 -1452 492 -1444
rect 191 -1456 388 -1454
rect 384 -1479 388 -1456
rect 450 -1461 456 -1452
rect 498 -1448 804 -1437
rect 498 -1473 505 -1448
rect 404 -1477 508 -1473
rect 176 -1493 202 -1492
rect 176 -1497 203 -1493
rect 176 -1498 182 -1497
rect 146 -1506 154 -1499
rect 195 -1500 203 -1497
rect 147 -1512 153 -1506
rect 195 -1531 202 -1500
rect 101 -1535 205 -1531
rect 384 -1532 387 -1479
rect 81 -1590 84 -1543
rect 81 -1594 92 -1590
rect 81 -1625 86 -1594
rect 92 -1613 98 -1602
rect 101 -1614 104 -1535
rect 167 -1544 184 -1543
rect 199 -1543 204 -1535
rect 384 -1536 395 -1532
rect 189 -1544 193 -1543
rect 167 -1547 193 -1544
rect 167 -1563 170 -1547
rect 107 -1568 170 -1563
rect 107 -1591 110 -1568
rect 141 -1590 144 -1574
rect 167 -1584 170 -1568
rect 132 -1594 144 -1590
rect 126 -1606 130 -1602
rect 108 -1610 130 -1606
rect 108 -1621 115 -1610
rect 126 -1613 130 -1610
rect 140 -1621 144 -1594
rect 81 -1647 84 -1625
rect 98 -1626 115 -1621
rect 132 -1625 144 -1621
rect 153 -1625 157 -1584
rect 163 -1587 170 -1584
rect 173 -1566 181 -1562
rect 163 -1599 166 -1587
rect 173 -1590 176 -1566
rect 181 -1585 187 -1574
rect 190 -1586 193 -1547
rect 196 -1547 251 -1543
rect 196 -1563 199 -1547
rect 221 -1566 233 -1562
rect 215 -1578 219 -1574
rect 197 -1582 219 -1578
rect 197 -1593 204 -1582
rect 215 -1585 219 -1582
rect 229 -1593 233 -1566
rect 187 -1598 204 -1593
rect 221 -1597 233 -1593
rect 163 -1603 170 -1599
rect 165 -1605 170 -1603
rect 81 -1651 92 -1647
rect 81 -1682 86 -1651
rect 92 -1670 98 -1659
rect 101 -1671 104 -1626
rect 107 -1648 110 -1626
rect 141 -1647 144 -1625
rect 132 -1651 144 -1647
rect 126 -1663 130 -1659
rect 108 -1667 130 -1663
rect 108 -1678 115 -1667
rect 126 -1670 130 -1667
rect 140 -1678 144 -1651
rect 148 -1629 158 -1625
rect 148 -1673 152 -1629
rect 158 -1648 164 -1637
rect 167 -1649 170 -1605
rect 198 -1609 201 -1598
rect 230 -1606 233 -1597
rect 173 -1614 245 -1609
rect 173 -1626 176 -1614
rect 222 -1621 233 -1617
rect 198 -1629 210 -1625
rect 192 -1641 196 -1637
rect 174 -1645 196 -1641
rect 174 -1656 181 -1645
rect 192 -1648 196 -1645
rect 206 -1656 210 -1629
rect 222 -1652 227 -1621
rect 233 -1640 239 -1629
rect 242 -1641 245 -1614
rect 248 -1618 251 -1547
rect 384 -1567 389 -1536
rect 395 -1555 401 -1544
rect 404 -1556 407 -1477
rect 470 -1486 487 -1485
rect 502 -1485 507 -1477
rect 492 -1486 496 -1485
rect 470 -1489 496 -1486
rect 470 -1505 473 -1489
rect 410 -1510 473 -1505
rect 410 -1533 413 -1510
rect 444 -1532 447 -1516
rect 470 -1526 473 -1510
rect 435 -1536 447 -1532
rect 429 -1548 433 -1544
rect 411 -1552 433 -1548
rect 411 -1563 418 -1552
rect 429 -1555 433 -1552
rect 443 -1563 447 -1536
rect 280 -1617 285 -1592
rect 273 -1621 285 -1617
rect 267 -1633 271 -1629
rect 249 -1637 271 -1633
rect 249 -1648 256 -1637
rect 267 -1640 271 -1637
rect 281 -1648 285 -1621
rect 384 -1589 387 -1567
rect 401 -1568 418 -1563
rect 435 -1567 447 -1563
rect 456 -1567 460 -1526
rect 466 -1529 473 -1526
rect 476 -1508 484 -1504
rect 466 -1541 469 -1529
rect 476 -1532 479 -1508
rect 484 -1527 490 -1516
rect 493 -1528 496 -1489
rect 499 -1489 554 -1485
rect 499 -1505 502 -1489
rect 524 -1508 536 -1504
rect 518 -1520 522 -1516
rect 500 -1524 522 -1520
rect 500 -1535 507 -1524
rect 518 -1527 522 -1524
rect 532 -1535 536 -1508
rect 490 -1540 507 -1535
rect 524 -1539 536 -1535
rect 466 -1545 473 -1541
rect 468 -1547 473 -1545
rect 384 -1593 395 -1589
rect 384 -1624 389 -1593
rect 395 -1612 401 -1601
rect 404 -1613 407 -1568
rect 410 -1590 413 -1568
rect 444 -1589 447 -1567
rect 435 -1593 447 -1589
rect 429 -1605 433 -1601
rect 411 -1609 433 -1605
rect 411 -1620 418 -1609
rect 429 -1612 433 -1609
rect 443 -1620 447 -1593
rect 451 -1571 461 -1567
rect 451 -1615 455 -1571
rect 461 -1590 467 -1579
rect 470 -1591 473 -1547
rect 501 -1551 504 -1540
rect 533 -1548 536 -1539
rect 476 -1556 548 -1551
rect 476 -1568 479 -1556
rect 525 -1563 536 -1559
rect 501 -1571 513 -1567
rect 495 -1583 499 -1579
rect 477 -1587 499 -1583
rect 477 -1598 484 -1587
rect 495 -1590 499 -1587
rect 509 -1598 513 -1571
rect 525 -1594 530 -1563
rect 536 -1582 542 -1571
rect 545 -1583 548 -1556
rect 551 -1560 554 -1489
rect 583 -1559 588 -1534
rect 576 -1563 588 -1559
rect 570 -1575 574 -1571
rect 552 -1579 574 -1575
rect 552 -1590 559 -1579
rect 570 -1582 574 -1579
rect 584 -1590 588 -1563
rect 542 -1595 559 -1590
rect 576 -1594 588 -1590
rect 467 -1603 484 -1598
rect 501 -1602 513 -1598
rect 451 -1620 465 -1615
rect 385 -1634 389 -1624
rect 401 -1625 418 -1620
rect 435 -1624 447 -1620
rect 239 -1653 256 -1648
rect 273 -1652 285 -1648
rect 164 -1661 181 -1656
rect 198 -1660 210 -1656
rect 148 -1678 162 -1673
rect 82 -1692 86 -1682
rect 98 -1683 115 -1678
rect 132 -1682 144 -1678
rect 19 -1702 87 -1692
rect 19 -1773 25 -1702
rect 104 -1714 111 -1683
rect 33 -1721 111 -1714
rect 157 -1710 163 -1678
rect 174 -1680 180 -1661
rect 207 -1669 210 -1660
rect 249 -1673 254 -1653
rect 282 -1662 285 -1652
rect 283 -1669 285 -1662
rect 218 -1679 254 -1673
rect 174 -1686 215 -1680
rect 192 -1695 203 -1691
rect 192 -1710 197 -1695
rect 157 -1716 197 -1710
rect 33 -1760 41 -1721
rect 192 -1726 197 -1716
rect 203 -1714 209 -1703
rect 212 -1715 215 -1686
rect 218 -1692 221 -1679
rect 243 -1695 255 -1691
rect 237 -1707 241 -1703
rect 219 -1711 241 -1707
rect 219 -1722 226 -1711
rect 237 -1714 241 -1711
rect 251 -1711 255 -1695
rect 282 -1711 285 -1669
rect 251 -1716 285 -1711
rect 251 -1722 255 -1716
rect 209 -1727 226 -1722
rect 243 -1726 255 -1722
rect 219 -1730 226 -1727
rect 106 -1737 226 -1730
rect 252 -1735 255 -1726
rect 80 -1749 90 -1740
rect 35 -1765 40 -1760
rect 85 -1761 90 -1749
rect 35 -1768 50 -1765
rect 19 -1776 31 -1773
rect 20 -1777 31 -1776
rect 20 -1808 25 -1777
rect 31 -1796 37 -1785
rect 40 -1797 43 -1768
rect 46 -1770 50 -1768
rect 46 -1774 49 -1770
rect 86 -1773 89 -1761
rect 71 -1777 83 -1773
rect 65 -1789 69 -1785
rect 47 -1793 69 -1789
rect 47 -1804 54 -1793
rect 65 -1796 69 -1793
rect 79 -1804 83 -1777
rect 20 -1833 23 -1808
rect 37 -1809 54 -1804
rect 71 -1808 83 -1804
rect 41 -1825 45 -1809
rect 79 -1820 83 -1808
rect 82 -1825 83 -1820
rect 86 -1777 97 -1773
rect 86 -1808 91 -1777
rect 97 -1796 103 -1785
rect 106 -1797 109 -1737
rect 112 -1751 180 -1748
rect 112 -1774 115 -1751
rect 172 -1755 180 -1751
rect 219 -1755 226 -1737
rect 146 -1758 149 -1757
rect 144 -1773 149 -1758
rect 172 -1759 198 -1755
rect 137 -1777 149 -1773
rect 172 -1775 175 -1759
rect 131 -1789 135 -1785
rect 113 -1793 135 -1789
rect 113 -1804 120 -1793
rect 131 -1796 135 -1793
rect 145 -1804 149 -1777
rect 7 -1837 23 -1833
rect 27 -1829 45 -1825
rect 7 -1854 11 -1837
rect 7 -1858 18 -1854
rect 7 -1886 12 -1858
rect 18 -1877 24 -1866
rect 27 -1878 30 -1829
rect 86 -1830 89 -1808
rect 103 -1809 120 -1804
rect 137 -1808 149 -1804
rect 33 -1837 81 -1833
rect 33 -1855 36 -1837
rect 58 -1858 70 -1854
rect 52 -1870 56 -1866
rect 34 -1874 56 -1870
rect 34 -1885 41 -1874
rect 52 -1877 56 -1874
rect 66 -1885 70 -1858
rect 7 -1899 14 -1886
rect 24 -1890 41 -1885
rect 58 -1889 70 -1885
rect 8 -1964 14 -1899
rect 67 -1898 70 -1889
rect 67 -1950 71 -1898
rect 74 -1940 81 -1837
rect 86 -1834 97 -1830
rect 86 -1912 91 -1834
rect 97 -1853 103 -1842
rect 106 -1854 109 -1809
rect 112 -1831 115 -1809
rect 146 -1830 149 -1808
rect 167 -1779 175 -1775
rect 178 -1778 186 -1774
rect 167 -1818 170 -1779
rect 178 -1809 181 -1778
rect 186 -1797 192 -1786
rect 195 -1798 198 -1759
rect 201 -1759 256 -1755
rect 282 -1759 285 -1716
rect 322 -1644 390 -1634
rect 322 -1715 328 -1644
rect 407 -1656 414 -1625
rect 336 -1663 414 -1656
rect 460 -1652 466 -1620
rect 477 -1622 483 -1603
rect 510 -1611 513 -1602
rect 552 -1615 557 -1595
rect 585 -1604 588 -1594
rect 586 -1611 588 -1604
rect 521 -1621 557 -1615
rect 477 -1628 518 -1622
rect 495 -1637 506 -1633
rect 495 -1652 500 -1637
rect 460 -1658 500 -1652
rect 336 -1702 344 -1663
rect 495 -1668 500 -1658
rect 506 -1656 512 -1645
rect 515 -1657 518 -1628
rect 521 -1634 524 -1621
rect 546 -1637 558 -1633
rect 540 -1649 544 -1645
rect 522 -1653 544 -1649
rect 522 -1664 529 -1653
rect 540 -1656 544 -1653
rect 554 -1653 558 -1637
rect 585 -1653 588 -1611
rect 554 -1658 588 -1653
rect 554 -1664 558 -1658
rect 512 -1669 529 -1664
rect 546 -1668 558 -1664
rect 522 -1672 529 -1669
rect 409 -1679 529 -1672
rect 555 -1677 558 -1668
rect 383 -1691 393 -1682
rect 338 -1707 343 -1702
rect 388 -1703 393 -1691
rect 338 -1710 353 -1707
rect 322 -1718 334 -1715
rect 201 -1775 204 -1759
rect 226 -1778 238 -1774
rect 220 -1790 224 -1786
rect 202 -1794 224 -1790
rect 202 -1805 209 -1794
rect 220 -1797 224 -1794
rect 234 -1805 238 -1778
rect 192 -1810 209 -1805
rect 226 -1809 238 -1805
rect 167 -1821 175 -1818
rect 203 -1821 206 -1810
rect 235 -1818 238 -1809
rect 247 -1821 250 -1814
rect 137 -1834 149 -1830
rect 131 -1846 135 -1842
rect 113 -1850 135 -1846
rect 113 -1861 120 -1850
rect 131 -1853 135 -1850
rect 145 -1861 149 -1834
rect 103 -1866 120 -1861
rect 137 -1865 149 -1861
rect 114 -1890 119 -1866
rect 152 -1841 163 -1837
rect 152 -1871 157 -1841
rect 163 -1860 169 -1849
rect 172 -1861 175 -1821
rect 178 -1826 250 -1821
rect 178 -1838 181 -1826
rect 227 -1833 238 -1829
rect 203 -1841 215 -1837
rect 197 -1853 201 -1849
rect 179 -1857 201 -1853
rect 179 -1868 186 -1857
rect 197 -1860 201 -1857
rect 211 -1868 215 -1841
rect 227 -1864 232 -1833
rect 238 -1852 244 -1841
rect 247 -1853 250 -1826
rect 253 -1830 256 -1759
rect 283 -1765 285 -1759
rect 282 -1800 285 -1765
rect 323 -1719 334 -1718
rect 323 -1750 328 -1719
rect 334 -1738 340 -1727
rect 343 -1739 346 -1710
rect 349 -1712 353 -1710
rect 349 -1716 352 -1712
rect 389 -1715 392 -1703
rect 374 -1719 386 -1715
rect 368 -1731 372 -1727
rect 350 -1735 372 -1731
rect 350 -1746 357 -1735
rect 368 -1738 372 -1735
rect 382 -1746 386 -1719
rect 323 -1775 326 -1750
rect 340 -1751 357 -1746
rect 374 -1750 386 -1746
rect 344 -1767 348 -1751
rect 382 -1762 386 -1750
rect 385 -1767 386 -1762
rect 389 -1719 400 -1715
rect 389 -1750 394 -1719
rect 400 -1738 406 -1727
rect 409 -1739 412 -1679
rect 415 -1693 483 -1690
rect 415 -1716 418 -1693
rect 475 -1697 483 -1693
rect 522 -1697 529 -1679
rect 449 -1700 452 -1699
rect 447 -1715 452 -1700
rect 475 -1701 501 -1697
rect 440 -1719 452 -1715
rect 475 -1717 478 -1701
rect 434 -1731 438 -1727
rect 416 -1735 438 -1731
rect 416 -1746 423 -1735
rect 434 -1738 438 -1735
rect 448 -1746 452 -1719
rect 310 -1779 326 -1775
rect 330 -1771 348 -1767
rect 310 -1796 314 -1779
rect 310 -1800 321 -1796
rect 282 -1804 290 -1800
rect 287 -1829 290 -1804
rect 278 -1833 290 -1829
rect 272 -1845 276 -1841
rect 254 -1849 276 -1845
rect 254 -1860 261 -1849
rect 272 -1852 276 -1849
rect 286 -1860 290 -1833
rect 310 -1828 315 -1800
rect 321 -1819 327 -1808
rect 330 -1820 333 -1771
rect 389 -1772 392 -1750
rect 406 -1751 423 -1746
rect 440 -1750 452 -1746
rect 336 -1779 384 -1775
rect 336 -1797 339 -1779
rect 361 -1800 373 -1796
rect 355 -1812 359 -1808
rect 337 -1816 359 -1812
rect 337 -1827 344 -1816
rect 355 -1819 359 -1816
rect 369 -1827 373 -1800
rect 310 -1841 317 -1828
rect 327 -1832 344 -1827
rect 361 -1831 373 -1827
rect 244 -1865 261 -1860
rect 278 -1864 290 -1860
rect 152 -1877 158 -1871
rect 169 -1873 186 -1868
rect 203 -1872 215 -1868
rect 152 -1881 174 -1877
rect 114 -1893 129 -1890
rect 99 -1902 110 -1898
rect 99 -1912 104 -1902
rect 86 -1916 104 -1912
rect 99 -1933 104 -1916
rect 110 -1921 116 -1910
rect 119 -1922 122 -1893
rect 125 -1895 129 -1893
rect 125 -1899 128 -1895
rect 150 -1902 162 -1898
rect 144 -1914 148 -1910
rect 126 -1918 148 -1914
rect 126 -1929 133 -1918
rect 144 -1921 148 -1918
rect 158 -1929 162 -1902
rect 116 -1934 133 -1929
rect 150 -1933 162 -1929
rect 122 -1940 129 -1934
rect 74 -1946 129 -1940
rect 122 -1947 129 -1946
rect 159 -1950 162 -1933
rect 67 -1955 162 -1950
rect 168 -1964 174 -1881
rect 179 -1892 185 -1873
rect 212 -1881 215 -1872
rect 254 -1885 259 -1865
rect 287 -1873 290 -1864
rect 288 -1880 290 -1873
rect 223 -1891 259 -1885
rect 179 -1895 220 -1892
rect 184 -1898 220 -1895
rect 197 -1907 208 -1903
rect 197 -1938 202 -1907
rect 208 -1926 214 -1915
rect 217 -1927 220 -1898
rect 223 -1904 226 -1891
rect 287 -1903 290 -1880
rect 248 -1907 290 -1903
rect 256 -1908 290 -1907
rect 311 -1906 317 -1841
rect 370 -1840 373 -1831
rect 370 -1892 374 -1840
rect 377 -1882 384 -1779
rect 389 -1776 400 -1772
rect 389 -1854 394 -1776
rect 400 -1795 406 -1784
rect 409 -1796 412 -1751
rect 415 -1773 418 -1751
rect 449 -1772 452 -1750
rect 470 -1721 478 -1717
rect 481 -1720 489 -1716
rect 470 -1760 473 -1721
rect 481 -1751 484 -1720
rect 489 -1739 495 -1728
rect 498 -1740 501 -1701
rect 504 -1701 559 -1697
rect 585 -1701 588 -1658
rect 504 -1717 507 -1701
rect 529 -1720 541 -1716
rect 523 -1732 527 -1728
rect 505 -1736 527 -1732
rect 505 -1747 512 -1736
rect 523 -1739 527 -1736
rect 537 -1747 541 -1720
rect 495 -1752 512 -1747
rect 529 -1751 541 -1747
rect 470 -1763 478 -1760
rect 506 -1763 509 -1752
rect 538 -1760 541 -1751
rect 550 -1763 553 -1756
rect 440 -1776 452 -1772
rect 434 -1788 438 -1784
rect 416 -1792 438 -1788
rect 416 -1803 423 -1792
rect 434 -1795 438 -1792
rect 448 -1803 452 -1776
rect 406 -1808 423 -1803
rect 440 -1807 452 -1803
rect 417 -1832 422 -1808
rect 455 -1783 466 -1779
rect 455 -1813 460 -1783
rect 466 -1802 472 -1791
rect 475 -1803 478 -1763
rect 481 -1768 553 -1763
rect 481 -1780 484 -1768
rect 530 -1775 541 -1771
rect 506 -1783 518 -1779
rect 500 -1795 504 -1791
rect 482 -1799 504 -1795
rect 482 -1810 489 -1799
rect 500 -1802 504 -1799
rect 514 -1810 518 -1783
rect 530 -1806 535 -1775
rect 541 -1794 547 -1783
rect 550 -1795 553 -1768
rect 556 -1772 559 -1701
rect 586 -1707 588 -1701
rect 585 -1742 588 -1707
rect 585 -1746 593 -1742
rect 590 -1771 593 -1746
rect 581 -1775 593 -1771
rect 575 -1787 579 -1783
rect 557 -1791 579 -1787
rect 557 -1802 564 -1791
rect 575 -1794 579 -1791
rect 589 -1802 593 -1775
rect 547 -1807 564 -1802
rect 581 -1806 593 -1802
rect 455 -1819 461 -1813
rect 472 -1815 489 -1810
rect 506 -1814 518 -1810
rect 455 -1823 477 -1819
rect 417 -1835 432 -1832
rect 402 -1844 413 -1840
rect 402 -1854 407 -1844
rect 389 -1858 407 -1854
rect 402 -1875 407 -1858
rect 413 -1863 419 -1852
rect 422 -1864 425 -1835
rect 428 -1837 432 -1835
rect 428 -1841 431 -1837
rect 453 -1844 465 -1840
rect 447 -1856 451 -1852
rect 429 -1860 451 -1856
rect 429 -1871 436 -1860
rect 447 -1863 451 -1860
rect 461 -1871 465 -1844
rect 419 -1876 436 -1871
rect 453 -1875 465 -1871
rect 425 -1882 432 -1876
rect 377 -1888 432 -1882
rect 425 -1889 432 -1888
rect 462 -1892 465 -1875
rect 370 -1897 465 -1892
rect 471 -1906 477 -1823
rect 482 -1834 488 -1815
rect 515 -1823 518 -1814
rect 557 -1827 562 -1807
rect 590 -1815 593 -1806
rect 591 -1822 593 -1815
rect 526 -1833 562 -1827
rect 482 -1837 523 -1834
rect 487 -1840 523 -1837
rect 500 -1849 511 -1845
rect 500 -1880 505 -1849
rect 511 -1868 517 -1857
rect 520 -1869 523 -1840
rect 526 -1846 529 -1833
rect 590 -1845 593 -1822
rect 551 -1849 593 -1845
rect 559 -1850 593 -1849
rect 545 -1861 549 -1857
rect 527 -1865 549 -1861
rect 527 -1876 534 -1865
rect 545 -1868 549 -1865
rect 559 -1876 563 -1850
rect 500 -1906 506 -1880
rect 517 -1881 534 -1876
rect 551 -1880 563 -1876
rect 242 -1919 246 -1915
rect 224 -1923 246 -1919
rect 224 -1934 231 -1923
rect 242 -1926 246 -1923
rect 256 -1934 260 -1908
rect 311 -1914 506 -1906
rect 311 -1915 505 -1914
rect 350 -1929 507 -1921
rect 197 -1964 203 -1938
rect 214 -1939 231 -1934
rect 248 -1938 260 -1934
rect 8 -1971 203 -1964
rect 18 -1972 203 -1971
rect 18 -1973 202 -1972
rect 47 -1987 204 -1979
rect 197 -1991 204 -1987
rect 196 -2014 204 -1991
rect -22 -2017 204 -2014
rect 217 -2013 223 -1939
rect 257 -1947 260 -1938
rect 500 -1950 507 -1929
rect 381 -1951 507 -1950
rect 372 -1955 507 -1951
rect 520 -1953 526 -1881
rect 560 -1889 563 -1880
rect 217 -2017 366 -2013
rect -22 -2019 197 -2017
rect -17 -2020 123 -2019
rect 360 -2024 366 -2017
rect -35 -2031 63 -2030
rect -35 -2034 174 -2031
rect 166 -2209 174 -2034
rect 360 -2068 365 -2024
rect 239 -2074 365 -2068
rect 372 -2061 378 -1955
rect 520 -1958 594 -1953
rect 446 -2030 490 -2027
rect 446 -2031 481 -2030
rect 446 -2039 450 -2031
rect 477 -2039 481 -2031
rect 458 -2045 469 -2041
rect 462 -2056 466 -2045
rect 462 -2058 482 -2056
rect 372 -2064 447 -2061
rect 462 -2063 508 -2058
rect 239 -2147 245 -2074
rect 254 -2083 321 -2081
rect 327 -2083 362 -2081
rect 254 -2084 362 -2083
rect 254 -2085 289 -2084
rect 254 -2093 258 -2085
rect 285 -2093 289 -2085
rect 266 -2099 277 -2095
rect 269 -2110 273 -2099
rect 311 -2085 346 -2084
rect 311 -2093 315 -2085
rect 342 -2093 346 -2085
rect 323 -2099 334 -2095
rect 326 -2110 330 -2099
rect 253 -2115 273 -2110
rect 254 -2117 273 -2115
rect 254 -2121 258 -2117
rect 310 -2115 330 -2110
rect 372 -2112 376 -2064
rect 438 -2070 470 -2067
rect 391 -2082 435 -2079
rect 391 -2083 426 -2082
rect 391 -2091 395 -2083
rect 422 -2091 426 -2083
rect 403 -2097 414 -2093
rect 407 -2108 411 -2097
rect 407 -2111 427 -2108
rect 438 -2111 443 -2070
rect 477 -2073 482 -2063
rect 458 -2079 469 -2073
rect 446 -2085 450 -2079
rect 446 -2090 481 -2085
rect 502 -2091 508 -2063
rect 520 -2060 564 -2057
rect 520 -2061 555 -2060
rect 520 -2069 524 -2061
rect 551 -2069 555 -2061
rect 532 -2075 543 -2071
rect 536 -2086 540 -2075
rect 502 -2094 521 -2091
rect 536 -2093 556 -2086
rect 509 -2100 544 -2097
rect 353 -2113 376 -2112
rect 288 -2117 330 -2115
rect 288 -2118 315 -2117
rect 353 -2115 392 -2113
rect 345 -2116 392 -2115
rect 407 -2114 443 -2111
rect 407 -2115 427 -2114
rect 345 -2118 356 -2116
rect 253 -2127 258 -2121
rect 310 -2121 315 -2118
rect 265 -2124 315 -2121
rect 372 -2121 415 -2119
rect 322 -2122 415 -2121
rect 322 -2124 376 -2122
rect 310 -2127 315 -2124
rect 266 -2133 277 -2127
rect 323 -2133 334 -2127
rect 285 -2139 289 -2133
rect 342 -2139 346 -2133
rect 254 -2141 289 -2139
rect 311 -2141 346 -2139
rect 254 -2144 362 -2141
rect 372 -2142 376 -2124
rect 422 -2125 427 -2115
rect 403 -2131 414 -2125
rect 391 -2136 395 -2131
rect 391 -2139 425 -2136
rect 438 -2136 443 -2114
rect 454 -2105 498 -2102
rect 454 -2106 489 -2105
rect 454 -2114 458 -2106
rect 485 -2114 489 -2106
rect 466 -2120 477 -2116
rect 470 -2131 474 -2120
rect 470 -2132 490 -2131
rect 509 -2132 515 -2100
rect 551 -2103 556 -2093
rect 438 -2139 455 -2136
rect 470 -2138 515 -2132
rect 532 -2109 543 -2103
rect 520 -2115 524 -2109
rect 520 -2120 555 -2115
rect 372 -2145 478 -2142
rect 372 -2147 378 -2145
rect 239 -2152 378 -2147
rect 485 -2148 490 -2138
rect 466 -2154 477 -2148
rect 454 -2160 458 -2154
rect 520 -2159 526 -2120
rect 488 -2160 526 -2159
rect 454 -2165 526 -2160
rect 294 -2209 300 -2175
rect 166 -2212 300 -2209
rect 497 -2178 508 -2171
rect 167 -2213 294 -2212
rect 497 -2293 502 -2178
rect 587 -2289 593 -1958
rect 817 -2269 823 -1358
rect 857 -1366 860 -1357
rect 816 -2296 824 -2269
rect 917 -2289 920 -763
rect 993 -2286 996 -557
<< m2contact >>
rect 137 -158 154 -149
rect 690 -162 707 -148
rect 918 -158 928 -147
rect 1001 -150 1010 -143
rect -265 -184 -250 -171
rect 212 -181 223 -172
rect 526 -188 546 -172
rect 817 -186 833 -171
rect -341 -208 -330 -201
rect -108 -209 -99 -201
rect -17 -209 -8 -201
rect 612 -203 622 -193
rect -493 -230 -478 -220
rect -415 -226 -404 -219
rect -187 -230 -174 -220
rect 53 -223 65 -211
rect -513 -324 -501 -313
rect -360 -323 -348 -314
rect -286 -321 -271 -314
rect 118 -324 130 -314
rect -437 -349 -422 -341
rect -132 -348 -119 -340
rect 192 -350 203 -341
rect 666 -352 684 -340
rect -206 -372 -193 -363
rect -38 -371 -27 -362
rect 507 -372 518 -363
rect 897 -370 906 -363
rect 37 -398 49 -388
rect 984 -389 993 -382
rect 586 -399 598 -390
rect 800 -396 809 -389
rect -510 -455 -501 -448
rect -489 -451 -481 -444
rect -434 -455 -425 -448
rect -413 -451 -405 -444
rect -359 -455 -350 -448
rect -338 -451 -330 -444
rect -526 -576 -517 -568
rect -282 -455 -273 -448
rect -261 -451 -253 -444
rect -450 -576 -441 -568
rect -375 -576 -366 -568
rect -205 -455 -196 -448
rect -184 -451 -176 -444
rect -129 -455 -120 -448
rect -108 -451 -100 -444
rect -298 -576 -289 -568
rect -506 -693 -497 -685
rect -221 -576 -212 -568
rect -145 -576 -136 -568
rect -38 -455 -29 -448
rect -17 -451 -9 -444
rect 42 -454 51 -447
rect 63 -450 71 -443
rect 121 -453 130 -446
rect 142 -449 150 -442
rect -54 -576 -45 -568
rect 197 -452 206 -445
rect 218 -448 226 -441
rect 26 -575 35 -567
rect 105 -574 114 -566
rect 181 -573 190 -565
rect 511 -451 520 -444
rect 532 -447 540 -440
rect 593 -451 602 -444
rect 614 -447 622 -440
rect 673 -451 682 -444
rect 694 -447 702 -440
rect 495 -572 504 -564
rect 577 -572 586 -564
rect 657 -572 666 -564
rect 802 -452 811 -445
rect 823 -448 831 -441
rect 899 -452 908 -445
rect 920 -448 928 -441
rect 984 -452 992 -446
rect 1002 -450 1007 -443
rect 786 -573 795 -565
rect 1243 -460 1272 -441
rect 883 -573 892 -565
rect -198 -904 -189 -896
rect 967 -575 976 -567
rect 135 -923 144 -915
rect 678 -962 687 -954
rect -17 -1279 -6 -1269
rect 76 -1395 91 -1387
rect -262 -1476 -253 -1468
rect -567 -1589 -558 -1581
rect 78 -1543 87 -1535
<< metal2 >>
rect -509 -433 -504 -324
rect -488 -425 -482 -230
rect -508 -448 -505 -433
rect -490 -437 -482 -425
rect -433 -427 -427 -349
rect -432 -431 -426 -427
rect -487 -444 -484 -437
rect -432 -448 -429 -431
rect -411 -434 -407 -226
rect -357 -431 -351 -323
rect -336 -428 -332 -208
rect -280 -426 -274 -321
rect -259 -426 -255 -184
rect -414 -437 -405 -434
rect -411 -444 -408 -437
rect -357 -448 -354 -431
rect -336 -432 -333 -428
rect -280 -431 -275 -426
rect -336 -434 -332 -432
rect -339 -437 -330 -434
rect -336 -444 -333 -437
rect -280 -448 -277 -431
rect -259 -432 -256 -426
rect -203 -431 -198 -372
rect -259 -434 -255 -432
rect -262 -437 -253 -434
rect -259 -444 -256 -437
rect -203 -448 -200 -431
rect -182 -432 -179 -230
rect -182 -434 -178 -432
rect -185 -437 -176 -434
rect -182 -444 -179 -437
rect -127 -448 -124 -348
rect -106 -432 -103 -209
rect -106 -434 -102 -432
rect -109 -437 -100 -434
rect -106 -444 -103 -437
rect -36 -448 -33 -371
rect -14 -431 -11 -209
rect -15 -434 -11 -431
rect -18 -437 -9 -434
rect -15 -444 -12 -437
rect 44 -447 47 -398
rect 65 -433 69 -211
rect 62 -436 71 -433
rect 65 -443 68 -436
rect 123 -446 126 -324
rect 144 -427 147 -158
rect 141 -435 150 -427
rect 144 -442 147 -435
rect 199 -445 202 -350
rect 220 -426 223 -181
rect 217 -434 226 -426
rect 220 -441 223 -434
rect 513 -444 516 -372
rect 533 -433 538 -188
rect 534 -440 537 -433
rect 595 -444 598 -399
rect 616 -440 619 -203
rect 675 -430 679 -352
rect 675 -444 678 -430
rect 696 -440 699 -162
rect 804 -445 807 -396
rect 824 -416 828 -186
rect 825 -441 828 -416
rect 901 -445 904 -370
rect 922 -441 925 -158
rect 987 -446 992 -389
rect 1003 -443 1008 -150
rect 1251 -477 1263 -460
rect -527 -573 -526 -571
rect -530 -576 -526 -573
rect -452 -573 -450 -571
rect -517 -576 -450 -573
rect -376 -573 -375 -571
rect -441 -576 -375 -573
rect -299 -573 -298 -571
rect -366 -576 -298 -573
rect -222 -573 -221 -571
rect -289 -576 -221 -573
rect -146 -573 -145 -571
rect -212 -576 -145 -573
rect -55 -573 -54 -571
rect -136 -576 -54 -573
rect 24 -572 26 -570
rect 13 -573 26 -572
rect -45 -575 26 -573
rect 104 -571 105 -569
rect 93 -572 105 -571
rect 35 -574 105 -572
rect 180 -570 181 -568
rect 172 -571 181 -570
rect 114 -573 181 -571
rect 494 -569 495 -567
rect 248 -570 495 -569
rect 190 -572 495 -570
rect 576 -569 577 -567
rect 504 -572 577 -569
rect 656 -569 657 -567
rect 586 -572 657 -569
rect 733 -569 786 -568
rect 666 -572 786 -569
rect 190 -573 491 -572
rect 114 -574 177 -573
rect 35 -575 98 -574
rect -45 -576 18 -575
rect -464 -637 -459 -576
rect -505 -643 -459 -637
rect -401 -613 -395 -612
rect -401 -622 -280 -613
rect -401 -623 -359 -622
rect -503 -685 -499 -643
rect -437 -763 -432 -670
rect -401 -677 -395 -623
rect -400 -689 -395 -677
rect -315 -729 -305 -640
rect -344 -736 -299 -729
rect -425 -740 -412 -739
rect -425 -744 -413 -740
rect -425 -761 -422 -744
rect -411 -756 -408 -746
rect -411 -759 -368 -756
rect -436 -834 -432 -763
rect -371 -780 -368 -759
rect -366 -818 -310 -812
rect -522 -899 -514 -860
rect -447 -908 -442 -839
rect -437 -891 -432 -834
rect -427 -914 -306 -909
rect -340 -947 -308 -939
rect -429 -958 -411 -954
rect -429 -971 -425 -958
rect -518 -978 -504 -975
rect -429 -978 -364 -971
rect -518 -997 -513 -978
rect -429 -982 -425 -978
rect -367 -997 -364 -978
rect -367 -1001 -362 -997
rect -441 -1034 -436 -1020
rect -362 -1030 -304 -1023
rect -441 -1037 -421 -1034
rect -427 -1043 -421 -1037
rect -548 -1051 -547 -1050
rect -570 -1147 -564 -1132
rect -555 -1137 -547 -1051
rect -285 -1082 -280 -622
rect -217 -866 -213 -576
rect 40 -662 50 -654
rect 114 -660 140 -655
rect -179 -679 -59 -675
rect -179 -846 -175 -679
rect -76 -680 -59 -679
rect -65 -708 -59 -680
rect 40 -704 48 -662
rect -18 -715 -1 -709
rect 49 -729 60 -723
rect 105 -725 110 -661
rect 135 -680 140 -660
rect -154 -752 -138 -746
rect -154 -794 -149 -752
rect -24 -769 -1 -764
rect -154 -799 -86 -794
rect -24 -810 -18 -775
rect 41 -792 45 -770
rect 49 -792 55 -729
rect 41 -796 62 -792
rect 172 -802 179 -729
rect 129 -809 179 -802
rect -24 -816 -17 -810
rect 186 -816 194 -573
rect -24 -825 194 -816
rect 225 -837 230 -573
rect 614 -614 617 -572
rect 882 -570 883 -568
rect 795 -573 883 -570
rect 892 -573 967 -570
rect 976 -575 1202 -572
rect 442 -642 452 -634
rect 516 -640 542 -635
rect 337 -671 343 -655
rect 235 -676 343 -671
rect 235 -799 240 -676
rect 337 -688 343 -676
rect 442 -684 450 -642
rect 384 -695 401 -689
rect 451 -709 462 -703
rect 507 -705 512 -641
rect 537 -660 542 -640
rect 248 -732 264 -726
rect 248 -774 253 -732
rect 378 -749 401 -744
rect 248 -779 316 -774
rect 236 -803 240 -799
rect 378 -802 384 -755
rect 443 -772 447 -750
rect 451 -772 457 -709
rect 443 -776 464 -772
rect 574 -782 581 -709
rect 531 -789 581 -782
rect 614 -802 618 -614
rect 845 -616 855 -608
rect 919 -614 945 -609
rect 740 -662 746 -629
rect 845 -658 853 -616
rect 787 -669 804 -663
rect 854 -683 865 -677
rect 910 -679 915 -615
rect 940 -634 945 -614
rect 651 -706 667 -700
rect 651 -748 656 -706
rect 781 -723 804 -718
rect 651 -753 719 -748
rect 781 -776 787 -729
rect 846 -746 850 -724
rect 854 -746 860 -683
rect 846 -750 867 -746
rect 977 -756 984 -683
rect 934 -763 984 -756
rect 1053 -776 1057 -575
rect 780 -780 1057 -776
rect 236 -807 287 -803
rect 377 -806 618 -802
rect 236 -808 267 -807
rect 137 -846 231 -837
rect -179 -849 3 -846
rect -217 -867 -192 -866
rect -217 -873 -191 -867
rect -215 -875 -191 -873
rect -195 -896 -191 -875
rect -129 -974 -124 -881
rect -92 -900 -87 -881
rect -7 -940 3 -849
rect 137 -880 143 -846
rect 279 -870 287 -807
rect 279 -877 336 -870
rect 138 -915 142 -880
rect 326 -888 336 -877
rect 571 -888 580 -887
rect -36 -947 9 -940
rect -117 -951 -104 -950
rect -117 -955 -105 -951
rect -117 -972 -114 -955
rect -103 -967 -100 -957
rect -103 -970 -60 -967
rect -128 -1045 -124 -974
rect -63 -991 -60 -970
rect 204 -993 209 -900
rect 241 -919 246 -900
rect 326 -901 580 -888
rect 837 -896 843 -780
rect 1252 -874 1263 -477
rect 685 -897 843 -896
rect 326 -959 336 -901
rect 297 -966 342 -959
rect 216 -970 229 -969
rect 216 -974 228 -970
rect 216 -991 219 -974
rect 230 -986 233 -976
rect 230 -989 273 -986
rect -58 -1029 -2 -1023
rect -291 -1089 -280 -1082
rect -570 -1149 -526 -1147
rect -570 -1156 -432 -1149
rect -570 -1157 -526 -1156
rect -564 -1542 -561 -1157
rect -440 -1172 -432 -1156
rect -440 -1470 -431 -1172
rect -291 -1372 -286 -1089
rect -214 -1110 -206 -1071
rect -139 -1119 -134 -1050
rect -129 -1102 -124 -1045
rect 205 -1064 209 -993
rect 270 -1010 273 -989
rect 275 -1048 331 -1042
rect -119 -1125 2 -1120
rect 119 -1129 127 -1090
rect 194 -1138 199 -1069
rect 204 -1121 209 -1064
rect 214 -1144 335 -1139
rect -32 -1158 0 -1150
rect -121 -1169 -103 -1165
rect -121 -1182 -117 -1169
rect 301 -1177 333 -1169
rect -210 -1189 -196 -1186
rect -121 -1189 -56 -1182
rect -210 -1208 -205 -1189
rect -121 -1193 -117 -1189
rect -59 -1208 -56 -1189
rect 212 -1188 230 -1184
rect 212 -1201 216 -1188
rect 123 -1208 137 -1205
rect 212 -1208 277 -1201
rect -59 -1212 -54 -1208
rect 123 -1227 128 -1208
rect 212 -1212 216 -1208
rect -133 -1245 -128 -1231
rect 274 -1227 277 -1208
rect 274 -1231 279 -1227
rect -54 -1241 4 -1234
rect -133 -1248 -113 -1245
rect -119 -1254 -113 -1248
rect -240 -1262 -239 -1261
rect -247 -1348 -239 -1262
rect 200 -1264 205 -1250
rect 279 -1260 337 -1253
rect 200 -1267 220 -1264
rect -291 -1380 -95 -1372
rect -13 -1414 -8 -1279
rect 214 -1273 220 -1267
rect 93 -1281 94 -1280
rect 86 -1367 94 -1281
rect 571 -1346 580 -901
rect 681 -901 843 -897
rect 681 -954 685 -901
rect 816 -902 843 -901
rect 869 -883 1263 -874
rect 747 -1032 752 -939
rect 784 -958 789 -939
rect 869 -998 879 -883
rect 840 -1005 885 -998
rect 759 -1009 772 -1008
rect 759 -1013 771 -1009
rect 759 -1030 762 -1013
rect 773 -1025 776 -1015
rect 773 -1028 816 -1025
rect 748 -1103 752 -1032
rect 813 -1049 816 -1028
rect 818 -1087 874 -1081
rect 662 -1168 670 -1129
rect 737 -1177 742 -1108
rect 747 -1160 752 -1103
rect 757 -1183 878 -1178
rect 844 -1216 876 -1208
rect 755 -1227 773 -1223
rect 755 -1240 759 -1227
rect 666 -1247 680 -1244
rect 755 -1247 820 -1240
rect 666 -1266 671 -1247
rect 755 -1251 759 -1247
rect 817 -1266 820 -1247
rect 817 -1270 822 -1266
rect 743 -1303 748 -1289
rect 822 -1299 880 -1292
rect 743 -1306 763 -1303
rect 344 -1355 580 -1346
rect 343 -1356 580 -1355
rect -72 -1418 -8 -1414
rect -367 -1469 -262 -1468
rect -393 -1470 -262 -1469
rect -440 -1476 -262 -1470
rect -440 -1477 -279 -1476
rect -440 -1478 -326 -1477
rect -71 -1483 -61 -1418
rect -371 -1491 -61 -1483
rect -564 -1581 -560 -1542
rect -371 -1553 -365 -1491
rect -498 -1659 -493 -1566
rect -461 -1585 -456 -1566
rect -371 -1625 -366 -1553
rect -193 -1603 -188 -1510
rect -156 -1529 -151 -1510
rect -71 -1569 -61 -1491
rect 81 -1535 85 -1395
rect 255 -1471 262 -1408
rect 184 -1480 262 -1471
rect -100 -1576 -55 -1569
rect -181 -1580 -168 -1579
rect -181 -1584 -169 -1580
rect -181 -1601 -178 -1584
rect -167 -1596 -164 -1586
rect -167 -1599 -124 -1596
rect -405 -1632 -360 -1625
rect -486 -1636 -473 -1635
rect -486 -1640 -474 -1636
rect -486 -1657 -483 -1640
rect -472 -1652 -469 -1642
rect -472 -1655 -429 -1652
rect -497 -1730 -493 -1659
rect -432 -1676 -429 -1655
rect -192 -1674 -188 -1603
rect -127 -1620 -124 -1599
rect 147 -1613 152 -1520
rect 184 -1539 189 -1480
rect 343 -1498 350 -1356
rect 571 -1443 580 -1356
rect 757 -1312 763 -1306
rect 636 -1320 637 -1319
rect 629 -1406 637 -1320
rect 571 -1449 582 -1443
rect 269 -1503 351 -1498
rect 269 -1579 279 -1503
rect 450 -1555 455 -1469
rect 487 -1481 492 -1462
rect 572 -1521 582 -1449
rect 543 -1528 588 -1521
rect 462 -1532 475 -1531
rect 462 -1536 474 -1532
rect 462 -1553 465 -1536
rect 476 -1548 479 -1538
rect 476 -1551 519 -1548
rect 240 -1586 285 -1579
rect 159 -1590 172 -1589
rect 159 -1594 171 -1590
rect 159 -1611 162 -1594
rect 173 -1606 176 -1596
rect 173 -1609 216 -1606
rect -122 -1658 -66 -1652
rect -427 -1714 -371 -1708
rect -583 -1795 -575 -1756
rect -508 -1804 -503 -1735
rect -498 -1787 -493 -1730
rect -278 -1739 -270 -1700
rect -203 -1748 -198 -1679
rect -193 -1731 -188 -1674
rect 148 -1684 152 -1613
rect 213 -1630 216 -1609
rect 451 -1626 455 -1555
rect 516 -1572 519 -1551
rect 521 -1610 577 -1604
rect 218 -1668 274 -1662
rect 62 -1749 70 -1710
rect -183 -1754 -62 -1749
rect 137 -1758 142 -1689
rect 147 -1741 152 -1684
rect 365 -1691 373 -1652
rect 440 -1700 445 -1631
rect 450 -1683 455 -1626
rect 460 -1706 581 -1701
rect 547 -1739 579 -1731
rect 458 -1750 476 -1746
rect 157 -1764 278 -1759
rect 458 -1763 462 -1750
rect 369 -1770 383 -1767
rect 458 -1770 523 -1763
rect -96 -1787 -64 -1779
rect 369 -1789 374 -1770
rect 458 -1774 462 -1770
rect -185 -1798 -167 -1794
rect 244 -1797 276 -1789
rect 520 -1789 523 -1770
rect 520 -1793 525 -1789
rect -488 -1810 -367 -1805
rect -185 -1811 -181 -1798
rect 155 -1808 173 -1804
rect -274 -1818 -260 -1815
rect -185 -1818 -120 -1811
rect -401 -1843 -369 -1835
rect -274 -1837 -269 -1818
rect -185 -1822 -181 -1818
rect -123 -1837 -120 -1818
rect 155 -1821 159 -1808
rect 66 -1828 80 -1825
rect 155 -1828 220 -1821
rect -123 -1841 -118 -1837
rect 66 -1847 71 -1828
rect 155 -1832 159 -1828
rect -490 -1854 -472 -1850
rect 217 -1847 220 -1828
rect 446 -1826 451 -1812
rect 525 -1822 583 -1815
rect 446 -1829 466 -1826
rect 460 -1835 466 -1829
rect 339 -1843 340 -1842
rect 217 -1851 222 -1847
rect -490 -1867 -486 -1854
rect -579 -1874 -565 -1871
rect -490 -1874 -425 -1867
rect -579 -1893 -574 -1874
rect -490 -1878 -486 -1874
rect -428 -1893 -425 -1874
rect -197 -1874 -192 -1860
rect -118 -1870 -60 -1863
rect -197 -1877 -177 -1874
rect -183 -1883 -177 -1877
rect 143 -1884 148 -1870
rect 222 -1880 280 -1873
rect 143 -1887 163 -1884
rect -304 -1891 -303 -1890
rect -428 -1897 -423 -1893
rect -502 -1930 -497 -1916
rect -423 -1926 -365 -1919
rect -502 -1933 -482 -1930
rect -488 -1939 -482 -1933
rect -609 -1947 -608 -1946
rect -616 -2033 -608 -1947
rect -311 -1977 -303 -1891
rect 157 -1893 163 -1887
rect 36 -1901 37 -1900
rect 9 -1995 15 -1983
rect 29 -1987 37 -1901
rect 275 -1964 281 -1917
rect 332 -1929 340 -1843
rect 275 -1965 327 -1964
rect 275 -1971 328 -1965
rect 9 -2000 190 -1995
rect 183 -2182 190 -2000
rect 321 -2054 328 -1971
rect 426 -2031 436 -2023
rect 500 -2029 526 -2024
rect 321 -2077 327 -2054
rect 426 -2073 434 -2031
rect 368 -2084 385 -2078
rect 435 -2098 446 -2092
rect 491 -2094 496 -2030
rect 521 -2049 526 -2029
rect 232 -2121 248 -2115
rect 232 -2163 237 -2121
rect 362 -2138 385 -2133
rect 232 -2168 300 -2163
rect 362 -2182 368 -2144
rect 427 -2161 431 -2139
rect 435 -2161 441 -2098
rect 427 -2165 448 -2161
rect 558 -2171 565 -2098
rect 515 -2178 565 -2171
rect 182 -2187 368 -2182
<< m123contact >>
rect -437 -670 -431 -662
rect -500 -713 -495 -707
rect -400 -694 -395 -689
rect -315 -640 -304 -629
rect -411 -712 -406 -706
rect -351 -736 -344 -729
rect -413 -746 -408 -740
rect -304 -742 -299 -736
rect -449 -839 -441 -832
rect -427 -767 -422 -761
rect -368 -781 -362 -775
rect -374 -818 -366 -811
rect -310 -819 -301 -812
rect -523 -860 -513 -852
rect -514 -899 -504 -890
rect -437 -898 -432 -891
rect -447 -915 -440 -908
rect -435 -915 -427 -908
rect -306 -915 -301 -909
rect -346 -947 -340 -939
rect -308 -947 -302 -939
rect -411 -958 -406 -952
rect -508 -975 -502 -970
rect -430 -987 -425 -982
rect -518 -1004 -513 -997
rect -362 -1004 -357 -997
rect -441 -1020 -435 -1015
rect -369 -1030 -362 -1023
rect -304 -1030 -296 -1023
rect -555 -1051 -548 -1040
rect -426 -1048 -421 -1043
rect -573 -1132 -561 -1121
rect 122 -620 144 -606
rect 50 -662 60 -654
rect 104 -661 114 -653
rect -65 -675 -59 -669
rect -65 -714 -59 -708
rect -24 -715 -18 -709
rect -1 -714 5 -708
rect 39 -710 48 -704
rect 60 -729 70 -721
rect 133 -688 143 -680
rect -138 -752 -132 -746
rect -24 -775 -18 -769
rect -1 -770 5 -764
rect 39 -770 45 -765
rect -92 -806 -86 -799
rect 103 -733 113 -725
rect 170 -729 180 -721
rect 62 -796 68 -791
rect 122 -809 129 -802
rect 452 -642 462 -634
rect 506 -641 516 -633
rect 337 -655 343 -649
rect 337 -694 343 -688
rect 378 -695 384 -689
rect 401 -694 407 -688
rect 441 -690 450 -684
rect 462 -709 472 -701
rect 535 -668 545 -660
rect 264 -732 270 -726
rect 378 -755 384 -749
rect 401 -750 407 -744
rect 441 -750 447 -745
rect 310 -786 316 -779
rect 505 -713 515 -705
rect 572 -709 582 -701
rect 464 -776 470 -771
rect 524 -789 531 -782
rect 855 -616 865 -608
rect 909 -615 919 -607
rect 740 -629 746 -623
rect 740 -668 746 -662
rect 781 -669 787 -663
rect 804 -668 810 -662
rect 844 -664 853 -658
rect 865 -683 875 -675
rect 938 -642 948 -634
rect 667 -706 673 -700
rect 781 -729 787 -723
rect 804 -724 810 -718
rect 844 -724 850 -719
rect 713 -760 719 -753
rect 908 -687 918 -679
rect 975 -683 985 -675
rect 867 -750 873 -745
rect 927 -763 934 -756
rect -129 -881 -123 -873
rect -92 -881 -87 -871
rect -192 -924 -187 -918
rect -92 -905 -87 -900
rect -103 -923 -98 -917
rect 204 -900 210 -892
rect 241 -900 246 -890
rect -43 -947 -36 -940
rect 141 -943 146 -937
rect -105 -957 -100 -951
rect 4 -953 9 -947
rect -141 -1050 -133 -1043
rect -119 -978 -114 -972
rect -60 -992 -54 -986
rect 241 -924 246 -919
rect 230 -942 235 -936
rect 290 -966 297 -959
rect 228 -976 233 -970
rect 337 -972 342 -966
rect -66 -1029 -58 -1022
rect -2 -1030 7 -1023
rect -215 -1071 -205 -1063
rect -547 -1137 -537 -1129
rect -206 -1110 -196 -1101
rect 192 -1069 200 -1062
rect 214 -997 219 -991
rect 273 -1011 279 -1005
rect 267 -1048 275 -1041
rect 331 -1049 340 -1042
rect 118 -1090 128 -1082
rect -129 -1109 -124 -1102
rect -139 -1126 -132 -1119
rect -127 -1126 -119 -1119
rect 2 -1126 7 -1120
rect 127 -1129 137 -1120
rect 204 -1128 209 -1121
rect 194 -1145 201 -1138
rect 206 -1145 214 -1138
rect 335 -1145 340 -1139
rect -38 -1158 -32 -1150
rect 0 -1158 6 -1150
rect -103 -1169 -98 -1163
rect -200 -1186 -194 -1181
rect 295 -1177 301 -1169
rect 333 -1177 339 -1169
rect -122 -1198 -117 -1193
rect -210 -1215 -205 -1208
rect 230 -1188 235 -1182
rect 133 -1205 139 -1200
rect -54 -1215 -49 -1208
rect -133 -1231 -127 -1226
rect 211 -1217 216 -1212
rect 123 -1234 128 -1227
rect 279 -1234 284 -1227
rect -61 -1241 -54 -1234
rect 4 -1241 12 -1234
rect -247 -1262 -240 -1251
rect -118 -1259 -113 -1254
rect 200 -1250 206 -1245
rect 272 -1260 279 -1253
rect 337 -1260 345 -1253
rect -239 -1348 -229 -1340
rect -95 -1379 -80 -1363
rect 86 -1281 93 -1270
rect 215 -1278 220 -1273
rect 747 -939 753 -931
rect 784 -939 789 -929
rect 684 -982 689 -976
rect 784 -963 789 -958
rect 773 -981 778 -975
rect 833 -1005 840 -998
rect 771 -1015 776 -1009
rect 880 -1011 885 -1005
rect 735 -1108 743 -1101
rect 757 -1036 762 -1030
rect 816 -1050 822 -1044
rect 810 -1087 818 -1080
rect 874 -1088 883 -1081
rect 661 -1129 671 -1121
rect 670 -1168 680 -1159
rect 747 -1167 752 -1160
rect 737 -1184 744 -1177
rect 749 -1184 757 -1177
rect 878 -1184 883 -1178
rect 838 -1216 844 -1208
rect 876 -1216 882 -1208
rect 773 -1227 778 -1221
rect 676 -1244 682 -1239
rect 754 -1256 759 -1251
rect 666 -1273 671 -1266
rect 822 -1273 827 -1266
rect 743 -1289 749 -1284
rect 815 -1299 822 -1292
rect 880 -1299 888 -1292
rect 94 -1367 104 -1359
rect -193 -1510 -187 -1502
rect -156 -1510 -151 -1500
rect -256 -1553 -251 -1547
rect -498 -1566 -492 -1558
rect -461 -1566 -456 -1556
rect -561 -1609 -556 -1603
rect -461 -1590 -456 -1585
rect -472 -1608 -467 -1602
rect -156 -1534 -151 -1529
rect -167 -1552 -162 -1546
rect 252 -1408 264 -1393
rect 147 -1520 153 -1512
rect 84 -1563 89 -1557
rect -107 -1576 -100 -1569
rect -169 -1586 -164 -1580
rect -60 -1582 -55 -1576
rect -412 -1632 -405 -1625
rect -474 -1642 -469 -1636
rect -365 -1638 -360 -1632
rect -510 -1735 -502 -1728
rect -488 -1663 -483 -1657
rect -429 -1677 -423 -1671
rect -205 -1679 -197 -1672
rect -183 -1607 -178 -1601
rect 629 -1320 636 -1309
rect 758 -1317 763 -1312
rect 637 -1406 647 -1398
rect 448 -1452 461 -1443
rect 450 -1469 456 -1461
rect 487 -1462 492 -1452
rect 184 -1544 189 -1539
rect 173 -1562 178 -1556
rect 387 -1505 392 -1499
rect 487 -1486 492 -1481
rect 476 -1504 481 -1498
rect 536 -1528 543 -1521
rect 474 -1538 479 -1532
rect 583 -1534 588 -1528
rect 233 -1586 240 -1579
rect 171 -1596 176 -1590
rect 280 -1592 285 -1586
rect -124 -1621 -118 -1615
rect -130 -1658 -122 -1651
rect -66 -1659 -57 -1652
rect -279 -1700 -269 -1692
rect -435 -1714 -427 -1707
rect -371 -1715 -362 -1708
rect -584 -1756 -574 -1748
rect -575 -1795 -565 -1786
rect -270 -1739 -260 -1730
rect 135 -1689 143 -1682
rect 157 -1617 162 -1611
rect 216 -1631 222 -1625
rect 438 -1631 446 -1624
rect 460 -1559 465 -1553
rect 519 -1573 525 -1567
rect 513 -1610 521 -1603
rect 577 -1611 586 -1604
rect 364 -1652 374 -1644
rect 210 -1668 218 -1661
rect 274 -1669 283 -1662
rect 61 -1710 71 -1702
rect -193 -1738 -188 -1731
rect -203 -1755 -196 -1748
rect -191 -1755 -183 -1748
rect 70 -1749 80 -1740
rect -62 -1755 -57 -1749
rect 373 -1691 383 -1682
rect 450 -1690 455 -1683
rect 440 -1707 447 -1700
rect 452 -1707 460 -1700
rect 581 -1707 586 -1701
rect 541 -1739 547 -1731
rect 579 -1739 585 -1731
rect 147 -1748 152 -1741
rect 476 -1750 481 -1744
rect 137 -1765 144 -1758
rect 149 -1765 157 -1758
rect 278 -1765 283 -1759
rect 379 -1767 385 -1762
rect -102 -1787 -96 -1779
rect -64 -1787 -58 -1779
rect -498 -1794 -493 -1787
rect 457 -1779 462 -1774
rect -167 -1798 -162 -1792
rect 238 -1797 244 -1789
rect 276 -1797 282 -1789
rect 369 -1796 374 -1789
rect 525 -1796 530 -1789
rect -508 -1811 -501 -1804
rect -496 -1811 -488 -1804
rect -367 -1811 -362 -1805
rect -264 -1815 -258 -1810
rect 173 -1808 178 -1802
rect -407 -1843 -401 -1835
rect -369 -1843 -363 -1835
rect -186 -1827 -181 -1822
rect -274 -1844 -269 -1837
rect 76 -1825 82 -1820
rect 446 -1812 452 -1807
rect -118 -1844 -113 -1837
rect 154 -1837 159 -1832
rect -472 -1854 -467 -1848
rect 66 -1854 71 -1847
rect 518 -1822 525 -1815
rect 583 -1822 591 -1815
rect 332 -1843 339 -1832
rect 461 -1840 466 -1835
rect 222 -1854 227 -1847
rect -569 -1871 -563 -1866
rect -197 -1860 -191 -1855
rect -491 -1883 -486 -1878
rect -579 -1900 -574 -1893
rect -125 -1870 -118 -1863
rect -60 -1870 -52 -1863
rect 143 -1870 149 -1865
rect -311 -1891 -304 -1880
rect -182 -1888 -177 -1883
rect 215 -1880 222 -1873
rect 280 -1880 288 -1873
rect -423 -1900 -418 -1893
rect -502 -1916 -496 -1911
rect -430 -1926 -423 -1919
rect -365 -1926 -357 -1919
rect -616 -1947 -609 -1936
rect -487 -1944 -482 -1939
rect 29 -1901 36 -1890
rect 158 -1898 163 -1893
rect -303 -1977 -293 -1969
rect 8 -1983 18 -1971
rect 272 -1917 285 -1908
rect 340 -1929 350 -1921
rect 37 -1987 47 -1979
rect -608 -2033 -598 -2025
rect 436 -2031 446 -2023
rect 490 -2030 500 -2022
rect 321 -2083 327 -2077
rect 362 -2084 368 -2078
rect 385 -2083 391 -2077
rect 425 -2079 434 -2073
rect 446 -2098 456 -2090
rect 519 -2057 529 -2049
rect 248 -2121 254 -2115
rect 362 -2144 368 -2138
rect 385 -2139 391 -2133
rect 425 -2139 431 -2134
rect 294 -2175 300 -2168
rect 489 -2102 499 -2094
rect 556 -2098 566 -2090
rect 448 -2165 454 -2160
rect 508 -2178 515 -2171
<< metal3 >>
rect 129 -632 138 -620
rect 198 -632 206 -631
rect 129 -642 206 -632
rect 138 -645 206 -642
rect -495 -712 -411 -708
rect 198 -813 206 -645
rect 198 -828 358 -813
rect 200 -829 358 -828
rect 349 -912 358 -829
rect -187 -923 -103 -919
rect 349 -926 460 -912
rect 146 -942 230 -938
rect 452 -1402 460 -926
rect 689 -981 773 -977
rect 451 -1407 460 -1402
rect 451 -1443 456 -1407
rect 392 -1504 476 -1500
rect -251 -1552 -167 -1548
rect 89 -1562 173 -1558
rect -556 -1608 -472 -1604
<< labels >>
flabel metal1 1402 -440 1405 -438 1 FreeSans 89 0 0 0 VDD
flabel metal1 910 -602 911 -600 1 FreeSans 89 0 0 0 W15
flabel metal1 813 -596 814 -594 1 FreeSans 89 0 0 0 w14
flabel metal1 684 -622 685 -620 1 FreeSans 89 0 0 0 W13
flabel metal1 604 -606 605 -605 1 FreeSans 89 0 0 0 W12
flabel metal1 522 -601 523 -599 1 FreeSans 89 0 0 0 W11
flabel metal1 514 -854 517 -851 1 FreeSans 89 0 0 0 S1
flabel metal1 312 -856 315 -853 1 FreeSans 89 0 0 0 C2
flabel metal1 714 -834 715 -833 1 FreeSans 89 0 0 0 C1
flabel metal2 1195 -575 1196 -574 1 FreeSans 89 0 0 0 GND
flabel metal1 207 -611 208 -610 1 FreeSans 89 0 0 0 W10
flabel metal1 -27 -612 -25 -610 1 FreeSans 89 0 0 0 W7
flabel metal1 52 -617 54 -615 1 FreeSans 89 0 0 0 W8
flabel metal1 110 -808 112 -806 1 FreeSans 89 0 0 0 S2
flabel metal1 -90 -819 -89 -818 1 FreeSans 89 0 0 0 C3
flabel metal1 257 -1392 258 -1391 1 FreeSans 89 0 0 0 C5
flabel metal1 277 -1433 278 -1432 1 FreeSans 89 0 0 0 S3
flabel metal1 131 -607 133 -605 1 FreeSans 89 0 0 0 W9
flabel metal1 -118 -606 -117 -604 1 FreeSans 89 0 0 0 W6
flabel metal1 -194 -607 -193 -605 1 FreeSans 89 0 0 0 W5
flabel metal1 503 -1954 504 -1953 1 FreeSans 89 0 0 0 C7
flabel metal1 -272 -607 -271 -606 1 FreeSans 89 0 0 0 W4
flabel metal1 -76 -1373 -75 -1372 1 FreeSans 89 0 0 0 C6
flabel metal1 -57 -1374 -56 -1373 1 FreeSans 89 0 0 0 S4
flabel metal1 200 -2012 201 -2011 1 FreeSans 89 0 0 0 C8
flabel metal1 219 -2013 220 -2012 1 FreeSans 89 0 0 0 S5
flabel metal1 295 -2211 296 -2210 1 FreeSans 89 0 0 0 C10
flabel metal1 -852 -149 -851 -147 1 FreeSans 89 0 0 0 A0
flabel metal1 -768 -362 -767 -360 1 FreeSans 89 0 0 0 B1
flabel metal1 -767 -387 -766 -385 1 FreeSans 89 0 0 0 B0
flabel metal1 -765 -339 -762 -336 1 FreeSans 89 0 0 0 B2
flabel metal1 -846 -171 -842 -168 1 FreeSans 89 0 0 0 A1
flabel metal1 -835 -200 -830 -195 1 FreeSans 89 0 0 0 A2
flabel metal1 -763 -312 -761 -310 1 FreeSans 89 0 0 0 B3
flabel metal1 -854 -218 -850 -214 1 FreeSans 89 0 0 0 A3
flabel metal1 -348 -607 -347 -606 1 FreeSans 89 0 0 0 W3
flabel metal1 -423 -593 -422 -592 1 FreeSans 89 0 0 0 W2
flabel metal1 -384 -1162 -383 -1161 1 FreeSans 89 0 0 0 C9
flabel metal1 -365 -1207 -364 -1206 1 FreeSans 89 0 0 0 S6
flabel metal1 800 -1431 801 -1430 1 FreeSans 89 0 0 0 C4
flabel metal1 -145 -2013 -143 -2012 1 FreeSans 89 0 0 0 C11
flabel metal1 -499 -624 -498 -623 1 FreeSans 89 0 0 0 W1
flabel metal1 817 -2295 818 -2294 1 FreeSans 89 0 0 0 p2
flabel metal1 994 -2285 995 -2283 1 FreeSans 89 0 0 0 P0
flabel metal1 918 -2287 919 -2286 1 FreeSans 89 0 0 0 P1
flabel metal1 499 -2291 500 -2289 1 FreeSans 89 0 0 0 P4
flabel metal1 590 -2287 591 -2286 1 FreeSans 89 0 0 0 P3
flabel metal1 -121 -2274 -119 -2273 1 FreeSans 89 0 0 0 P5
flabel metal1 -427 -2260 -424 -2257 1 FreeSans 89 0 0 0 P6
flabel metal1 -445 -2260 -442 -2257 1 FreeSans 89 0 0 0 P7
<< end >>
